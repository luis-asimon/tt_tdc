VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_lcasimon_Tdc
  CLASS BLOCK ;
  FOREIGN tt_um_lcasimon_Tdc ;
  ORIGIN -1.000 0.100 ;
  SIZE 157.900 BY 226.470 ;
  OBS
      LAYER pwell ;
        RECT 107.460 173.770 110.295 174.200 ;
        RECT 107.460 169.420 107.890 173.770 ;
        RECT 108.065 169.620 109.325 173.570 ;
        RECT 107.460 168.990 110.295 169.420 ;
      LAYER nwell ;
        RECT 110.395 168.940 114.355 174.250 ;
        RECT 56.000 113.690 62.890 151.850 ;
      LAYER pwell ;
        RECT 64.305 151.370 67.005 151.800 ;
        RECT 64.305 142.780 64.735 151.370 ;
        RECT 65.275 142.980 66.035 151.170 ;
        RECT 66.575 142.780 67.005 151.370 ;
        RECT 91.785 151.370 94.485 151.800 ;
        RECT 64.305 142.350 67.005 142.780 ;
        RECT 72.460 142.650 77.900 143.080 ;
        RECT 64.305 138.160 67.005 138.590 ;
        RECT 64.305 117.890 64.735 138.160 ;
        RECT 65.275 118.090 66.035 137.960 ;
        RECT 66.575 117.890 67.005 138.160 ;
        RECT 64.305 117.460 67.005 117.890 ;
      LAYER nwell ;
        RECT 68.010 117.410 71.310 138.640 ;
        RECT 56.000 111.820 67.465 113.690 ;
      LAYER pwell ;
        RECT 67.540 113.210 70.375 113.640 ;
      LAYER nwell ;
        RECT 63.505 89.020 67.465 111.820 ;
      LAYER pwell ;
        RECT 68.985 89.700 69.745 113.010 ;
        RECT 69.945 89.500 70.375 113.210 ;
        RECT 72.460 113.340 72.890 142.650 ;
        RECT 73.430 113.500 74.190 142.490 ;
        RECT 76.170 113.900 76.930 142.090 ;
        RECT 77.470 113.340 77.900 142.650 ;
        RECT 72.460 112.910 77.900 113.340 ;
        RECT 80.890 142.650 86.330 143.080 ;
        RECT 80.890 113.340 81.320 142.650 ;
        RECT 81.860 113.900 82.620 142.090 ;
        RECT 84.600 113.500 85.360 142.490 ;
        RECT 85.900 113.340 86.330 142.650 ;
        RECT 91.785 142.780 92.215 151.370 ;
        RECT 92.755 142.980 93.515 151.170 ;
        RECT 94.055 142.780 94.485 151.370 ;
        RECT 91.785 142.350 94.485 142.780 ;
      LAYER nwell ;
        RECT 87.480 117.410 90.780 138.640 ;
      LAYER pwell ;
        RECT 91.785 138.160 94.485 138.590 ;
        RECT 91.785 117.890 92.215 138.160 ;
        RECT 92.755 118.090 93.515 137.960 ;
        RECT 94.055 117.890 94.485 138.160 ;
        RECT 91.785 117.460 94.485 117.890 ;
      LAYER nwell ;
        RECT 95.900 113.690 102.790 151.850 ;
      LAYER pwell ;
        RECT 80.890 112.910 86.330 113.340 ;
        RECT 88.415 113.210 91.250 113.640 ;
        RECT 67.540 89.070 70.375 89.500 ;
        RECT 88.415 89.500 88.845 113.210 ;
        RECT 89.045 89.700 89.805 113.010 ;
      LAYER nwell ;
        RECT 91.325 111.820 102.790 113.690 ;
        RECT 108.455 113.875 114.195 165.100 ;
      LAYER pwell ;
        RECT 121.710 164.580 125.980 165.010 ;
        RECT 114.795 118.220 117.695 118.455 ;
        RECT 121.710 118.220 122.140 164.580 ;
        RECT 114.795 118.025 122.140 118.220 ;
        RECT 114.795 114.615 115.225 118.025 ;
        RECT 115.765 114.775 116.725 117.865 ;
        RECT 117.265 117.790 122.140 118.025 ;
        RECT 117.265 114.615 118.495 117.790 ;
        RECT 114.795 114.185 118.495 114.615 ;
        RECT 88.415 89.070 91.250 89.500 ;
      LAYER nwell ;
        RECT 91.325 89.020 95.285 111.820 ;
        RECT 108.455 109.425 117.745 113.875 ;
      LAYER pwell ;
        RECT 118.065 110.080 118.495 114.185 ;
        RECT 119.035 110.240 120.295 117.630 ;
        RECT 120.835 110.080 122.140 117.790 ;
        RECT 118.065 109.650 122.140 110.080 ;
        RECT 71.345 82.540 74.460 82.970 ;
        RECT 71.345 78.190 71.775 82.540 ;
        RECT 72.315 78.390 73.575 82.340 ;
        RECT 71.345 77.760 74.460 78.190 ;
      LAYER nwell ;
        RECT 74.680 77.710 83.880 83.020 ;
      LAYER pwell ;
        RECT 84.100 82.540 87.215 82.970 ;
        RECT 84.985 78.390 86.245 82.340 ;
        RECT 86.785 78.190 87.215 82.540 ;
        RECT 84.100 77.760 87.215 78.190 ;
        RECT 88.375 82.890 91.210 83.320 ;
        RECT 88.375 78.540 88.805 82.890 ;
        RECT 88.980 78.740 90.240 82.690 ;
        RECT 88.375 78.110 91.210 78.540 ;
      LAYER nwell ;
        RECT 91.310 78.060 95.270 83.370 ;
        RECT 108.455 79.675 114.195 109.425 ;
      LAYER pwell ;
        RECT 114.795 84.020 117.695 84.255 ;
        RECT 121.710 84.020 122.140 109.650 ;
        RECT 114.795 83.825 122.140 84.020 ;
        RECT 114.795 80.415 115.225 83.825 ;
        RECT 115.765 80.575 116.725 83.665 ;
        RECT 117.265 83.590 122.140 83.825 ;
        RECT 117.265 80.415 118.495 83.590 ;
        RECT 114.795 79.985 118.495 80.415 ;
        RECT 64.595 72.230 67.430 72.660 ;
        RECT 64.595 63.580 65.025 72.230 ;
        RECT 65.200 63.780 66.460 72.030 ;
        RECT 64.595 63.150 67.430 63.580 ;
      LAYER nwell ;
        RECT 67.530 63.100 71.490 72.710 ;
      LAYER pwell ;
        RECT 73.615 72.230 76.450 72.660 ;
        RECT 73.615 63.580 74.045 72.230 ;
        RECT 74.220 63.780 75.480 72.030 ;
        RECT 73.615 63.150 76.450 63.580 ;
      LAYER nwell ;
        RECT 76.550 63.100 83.940 72.710 ;
      LAYER pwell ;
        RECT 84.040 72.230 86.875 72.660 ;
        RECT 85.010 63.780 86.270 72.030 ;
        RECT 86.445 63.580 86.875 72.230 ;
        RECT 84.040 63.150 86.875 63.580 ;
        RECT 88.375 72.230 91.210 72.660 ;
        RECT 88.375 63.580 88.805 72.230 ;
        RECT 88.980 63.780 90.240 72.030 ;
        RECT 88.375 63.150 91.210 63.580 ;
      LAYER nwell ;
        RECT 91.310 63.100 95.270 72.710 ;
        RECT 108.455 70.700 117.745 79.675 ;
      LAYER pwell ;
        RECT 118.065 75.880 118.495 79.985 ;
        RECT 119.035 76.040 120.295 83.430 ;
        RECT 120.835 77.110 122.140 83.590 ;
        RECT 122.680 77.270 123.640 164.420 ;
        RECT 124.050 77.270 125.010 164.420 ;
        RECT 125.550 77.110 125.980 164.580 ;
        RECT 120.835 76.680 125.980 77.110 ;
        RECT 120.835 75.880 121.265 76.680 ;
        RECT 118.065 75.450 121.265 75.880 ;
      LAYER nwell ;
        RECT 108.455 65.390 124.005 70.700 ;
      LAYER pwell ;
        RECT 124.325 70.180 127.225 70.610 ;
      LAYER nwell ;
        RECT 108.455 62.910 117.745 65.390 ;
      LAYER pwell ;
        RECT 124.325 65.360 124.755 70.180 ;
      LAYER nwell ;
        RECT 114.590 59.990 117.745 62.910 ;
      LAYER pwell ;
        RECT 118.340 64.930 124.755 65.360 ;
        RECT 118.340 60.660 118.770 64.930 ;
        RECT 119.310 60.820 120.270 64.770 ;
        RECT 122.025 60.820 122.985 64.770 ;
        RECT 123.525 60.750 124.755 64.930 ;
        RECT 125.295 60.910 126.255 70.020 ;
        RECT 126.795 60.750 127.225 70.180 ;
        RECT 123.525 60.660 127.225 60.750 ;
        RECT 118.340 60.320 127.225 60.660 ;
        RECT 118.340 60.230 123.955 60.320 ;
      LAYER li1 ;
        RECT 107.590 173.900 110.165 174.070 ;
        RECT 110.575 173.900 114.175 174.070 ;
        RECT 107.590 169.290 107.760 173.900 ;
        RECT 108.195 173.230 109.195 173.400 ;
        RECT 111.545 173.230 113.545 173.400 ;
        RECT 108.195 172.800 109.195 172.970 ;
        RECT 109.365 172.620 109.695 173.150 ;
        RECT 111.045 172.620 111.375 173.150 ;
        RECT 111.545 172.800 113.545 172.970 ;
        RECT 108.195 172.370 109.195 172.540 ;
        RECT 111.545 172.370 113.545 172.540 ;
        RECT 108.195 171.940 109.195 172.110 ;
        RECT 109.365 171.760 109.695 172.290 ;
        RECT 111.045 171.760 111.375 172.290 ;
        RECT 111.545 171.940 113.545 172.110 ;
        RECT 108.195 171.510 109.195 171.680 ;
        RECT 111.545 171.510 113.545 171.680 ;
        RECT 108.195 171.080 109.195 171.250 ;
        RECT 109.365 170.900 109.695 171.430 ;
        RECT 111.045 170.900 111.375 171.430 ;
        RECT 111.545 171.080 113.545 171.250 ;
        RECT 108.195 170.650 109.195 170.820 ;
        RECT 111.545 170.650 113.545 170.820 ;
        RECT 108.195 170.220 109.195 170.390 ;
        RECT 109.365 170.040 109.695 170.570 ;
        RECT 111.045 170.040 111.375 170.570 ;
        RECT 111.545 170.220 113.545 170.390 ;
        RECT 108.195 169.790 109.195 169.960 ;
        RECT 111.545 169.790 113.545 169.960 ;
        RECT 114.005 169.290 114.175 173.900 ;
        RECT 107.590 169.120 110.165 169.290 ;
        RECT 110.575 169.120 114.175 169.290 ;
        RECT 108.635 164.750 114.015 164.920 ;
        RECT 56.180 151.500 62.710 151.670 ;
        RECT 56.180 112.170 56.350 151.500 ;
        RECT 60.740 150.830 61.740 151.000 ;
        RECT 60.240 149.690 60.570 150.580 ;
        RECT 60.740 150.050 61.740 150.220 ;
        RECT 60.740 149.270 61.740 149.440 ;
        RECT 61.910 147.410 62.240 149.020 ;
        RECT 60.740 146.990 61.740 147.160 ;
        RECT 61.910 145.130 62.240 146.740 ;
        RECT 60.740 144.710 61.740 144.880 ;
        RECT 60.240 143.570 60.570 144.460 ;
        RECT 60.740 143.930 61.740 144.100 ;
        RECT 60.740 143.150 61.740 143.320 ;
        RECT 60.240 142.010 60.570 142.900 ;
        RECT 60.740 142.370 61.740 142.540 ;
        RECT 57.150 141.590 58.150 141.760 ;
        RECT 60.740 141.590 61.740 141.760 ;
        RECT 58.320 139.730 58.650 141.340 ;
        RECT 60.240 139.730 60.570 141.340 ;
        RECT 61.910 139.730 62.240 141.340 ;
        RECT 57.150 139.310 58.150 139.480 ;
        RECT 60.740 139.310 61.740 139.480 ;
        RECT 58.320 137.450 58.650 139.060 ;
        RECT 60.240 137.450 60.570 139.060 ;
        RECT 61.910 137.450 62.240 139.060 ;
        RECT 57.150 137.030 58.150 137.200 ;
        RECT 60.740 137.030 61.740 137.200 ;
        RECT 58.320 135.170 58.650 136.780 ;
        RECT 60.240 135.170 60.570 136.780 ;
        RECT 61.910 135.170 62.240 136.780 ;
        RECT 57.150 134.750 58.150 134.920 ;
        RECT 60.740 134.750 61.740 134.920 ;
        RECT 58.320 132.890 58.650 134.500 ;
        RECT 60.240 132.890 60.570 134.500 ;
        RECT 61.910 132.890 62.240 134.500 ;
        RECT 57.150 132.470 58.150 132.640 ;
        RECT 60.740 132.470 61.740 132.640 ;
        RECT 58.320 130.610 58.650 132.220 ;
        RECT 60.240 130.610 60.570 132.220 ;
        RECT 61.910 130.610 62.240 132.220 ;
        RECT 57.150 130.190 58.150 130.360 ;
        RECT 60.740 130.190 61.740 130.360 ;
        RECT 56.650 128.330 56.980 129.940 ;
        RECT 60.240 128.330 60.570 129.940 ;
        RECT 61.910 128.330 62.240 129.940 ;
        RECT 57.150 127.910 58.150 128.080 ;
        RECT 60.740 127.910 61.740 128.080 ;
        RECT 56.650 126.050 56.980 127.660 ;
        RECT 60.240 126.050 60.570 127.660 ;
        RECT 61.910 126.050 62.240 127.660 ;
        RECT 57.150 125.630 58.150 125.800 ;
        RECT 60.740 125.630 61.740 125.800 ;
        RECT 58.320 123.770 58.650 125.380 ;
        RECT 60.240 123.770 60.570 125.380 ;
        RECT 61.910 123.770 62.240 125.380 ;
        RECT 57.150 123.350 58.150 123.520 ;
        RECT 60.740 123.350 61.740 123.520 ;
        RECT 58.320 121.490 58.650 123.100 ;
        RECT 60.240 121.490 60.570 123.100 ;
        RECT 61.910 121.490 62.240 123.100 ;
        RECT 57.150 121.070 58.150 121.240 ;
        RECT 60.740 121.070 61.740 121.240 ;
        RECT 58.320 119.210 58.650 120.820 ;
        RECT 60.240 119.210 60.570 120.820 ;
        RECT 61.910 119.210 62.240 120.820 ;
        RECT 57.150 118.790 58.150 118.960 ;
        RECT 60.740 118.790 61.740 118.960 ;
        RECT 58.320 116.930 58.650 118.540 ;
        RECT 60.240 116.930 60.570 118.540 ;
        RECT 61.910 116.930 62.240 118.540 ;
        RECT 57.150 116.510 58.150 116.680 ;
        RECT 60.740 116.510 61.740 116.680 ;
        RECT 58.320 114.650 58.650 116.260 ;
        RECT 60.240 114.650 60.570 116.260 ;
        RECT 61.910 114.650 62.240 116.260 ;
        RECT 57.150 114.230 58.150 114.400 ;
        RECT 60.740 114.230 61.740 114.400 ;
        RECT 60.240 113.090 60.570 113.980 ;
        RECT 60.740 113.450 61.740 113.620 ;
        RECT 60.740 112.670 61.740 112.840 ;
        RECT 62.540 112.170 62.710 151.500 ;
        RECT 64.435 151.500 66.875 151.670 ;
        RECT 64.435 142.650 64.605 151.500 ;
        RECT 65.405 150.830 65.905 151.000 ;
        RECT 65.405 150.050 65.905 150.220 ;
        RECT 66.075 149.690 66.405 150.580 ;
        RECT 65.405 149.270 65.905 149.440 ;
        RECT 64.905 147.410 65.235 149.020 ;
        RECT 65.405 146.990 65.905 147.160 ;
        RECT 64.905 145.130 65.235 146.740 ;
        RECT 65.405 144.710 65.905 144.880 ;
        RECT 65.405 143.930 65.905 144.100 ;
        RECT 66.075 143.570 66.405 144.460 ;
        RECT 65.405 143.150 65.905 143.320 ;
        RECT 66.705 142.650 66.875 151.500 ;
        RECT 91.915 151.500 94.355 151.670 ;
        RECT 64.435 142.480 66.875 142.650 ;
        RECT 72.590 142.780 77.770 142.950 ;
        RECT 64.435 138.290 66.875 138.460 ;
        RECT 64.435 117.760 64.605 138.290 ;
        RECT 65.405 137.620 65.905 137.790 ;
        RECT 64.905 135.435 65.235 137.405 ;
        RECT 65.405 136.340 65.905 136.510 ;
        RECT 66.075 135.435 66.405 137.405 ;
        RECT 65.405 135.060 65.905 135.230 ;
        RECT 64.905 133.200 65.235 134.810 ;
        RECT 66.075 133.200 66.405 134.810 ;
        RECT 65.405 132.780 65.905 132.950 ;
        RECT 64.905 130.920 65.235 132.530 ;
        RECT 66.075 130.920 66.405 132.530 ;
        RECT 65.405 130.500 65.905 130.670 ;
        RECT 64.905 128.315 65.235 130.285 ;
        RECT 65.405 129.220 65.905 129.390 ;
        RECT 66.075 128.315 66.405 130.285 ;
        RECT 65.405 127.940 65.905 128.110 ;
        RECT 64.905 125.755 65.235 127.725 ;
        RECT 65.405 126.660 65.905 126.830 ;
        RECT 66.075 125.755 66.405 127.725 ;
        RECT 65.405 125.380 65.905 125.550 ;
        RECT 64.905 123.520 65.235 125.130 ;
        RECT 65.405 123.100 65.905 123.270 ;
        RECT 64.905 121.240 65.235 122.850 ;
        RECT 65.405 120.820 65.905 120.990 ;
        RECT 64.905 118.635 65.235 120.605 ;
        RECT 65.405 119.540 65.905 119.710 ;
        RECT 66.075 118.635 66.405 120.605 ;
        RECT 65.405 118.260 65.905 118.430 ;
        RECT 66.705 117.760 66.875 138.290 ;
        RECT 64.435 117.590 66.875 117.760 ;
        RECT 68.190 138.290 71.130 138.460 ;
        RECT 68.190 117.760 68.360 138.290 ;
        RECT 69.160 137.620 70.160 137.790 ;
        RECT 68.660 135.435 68.990 137.405 ;
        RECT 69.160 136.340 70.160 136.510 ;
        RECT 70.330 135.435 70.660 137.405 ;
        RECT 69.160 135.060 70.160 135.230 ;
        RECT 68.660 133.200 68.990 134.810 ;
        RECT 70.330 133.200 70.660 134.810 ;
        RECT 69.160 132.780 70.160 132.950 ;
        RECT 68.660 130.920 68.990 132.530 ;
        RECT 70.330 130.920 70.660 132.530 ;
        RECT 69.160 130.500 70.160 130.670 ;
        RECT 68.660 128.315 68.990 130.285 ;
        RECT 69.160 129.220 70.160 129.390 ;
        RECT 70.330 128.315 70.660 130.285 ;
        RECT 69.160 127.940 70.160 128.110 ;
        RECT 68.660 125.755 68.990 127.725 ;
        RECT 69.160 126.660 70.160 126.830 ;
        RECT 70.330 125.755 70.660 127.725 ;
        RECT 69.160 125.380 70.160 125.550 ;
        RECT 70.330 123.520 70.660 125.130 ;
        RECT 69.160 123.100 70.160 123.270 ;
        RECT 70.330 121.240 70.660 122.850 ;
        RECT 69.160 120.820 70.160 120.990 ;
        RECT 68.660 118.635 68.990 120.605 ;
        RECT 69.160 119.540 70.160 119.710 ;
        RECT 70.330 118.635 70.660 120.605 ;
        RECT 69.160 118.260 70.160 118.430 ;
        RECT 70.960 117.760 71.130 138.290 ;
        RECT 68.190 117.590 71.130 117.760 ;
        RECT 56.180 112.000 62.710 112.170 ;
        RECT 63.685 113.340 67.285 113.510 ;
        RECT 67.670 113.340 70.245 113.510 ;
        RECT 63.685 89.370 63.855 113.340 ;
        RECT 64.315 112.670 65.315 112.840 ;
        RECT 69.115 112.670 69.615 112.840 ;
        RECT 65.485 110.810 65.815 112.420 ;
        RECT 68.615 110.810 68.945 112.420 ;
        RECT 64.315 110.390 65.315 110.560 ;
        RECT 69.115 110.390 69.615 110.560 ;
        RECT 65.485 108.530 65.815 110.140 ;
        RECT 68.615 108.530 68.945 110.140 ;
        RECT 64.315 108.110 65.315 108.280 ;
        RECT 69.115 108.110 69.615 108.280 ;
        RECT 65.485 106.250 65.815 107.860 ;
        RECT 68.615 106.250 68.945 107.860 ;
        RECT 64.315 105.830 65.315 106.000 ;
        RECT 69.115 105.830 69.615 106.000 ;
        RECT 65.485 103.970 65.815 105.580 ;
        RECT 68.615 103.970 68.945 105.580 ;
        RECT 64.315 103.550 65.315 103.720 ;
        RECT 69.115 103.550 69.615 103.720 ;
        RECT 65.485 101.690 65.815 103.300 ;
        RECT 68.615 101.690 68.945 103.300 ;
        RECT 64.315 101.270 65.315 101.440 ;
        RECT 69.115 101.270 69.615 101.440 ;
        RECT 65.485 99.410 65.815 101.020 ;
        RECT 68.615 99.410 68.945 101.020 ;
        RECT 64.315 98.990 65.315 99.160 ;
        RECT 69.115 98.990 69.615 99.160 ;
        RECT 65.485 97.130 65.815 98.740 ;
        RECT 68.615 97.130 68.945 98.740 ;
        RECT 64.315 96.710 65.315 96.880 ;
        RECT 69.115 96.710 69.615 96.880 ;
        RECT 65.485 94.850 65.815 96.460 ;
        RECT 68.615 94.850 68.945 96.460 ;
        RECT 64.315 94.430 65.315 94.600 ;
        RECT 69.115 94.430 69.615 94.600 ;
        RECT 65.485 92.570 65.815 94.180 ;
        RECT 68.615 92.570 68.945 94.180 ;
        RECT 64.315 92.150 65.315 92.320 ;
        RECT 69.115 92.150 69.615 92.320 ;
        RECT 65.485 90.290 65.815 91.900 ;
        RECT 68.615 90.290 68.945 91.900 ;
        RECT 64.315 89.870 65.315 90.040 ;
        RECT 69.115 89.870 69.615 90.040 ;
        RECT 70.075 89.370 70.245 113.340 ;
        RECT 72.590 113.210 72.760 142.780 ;
        RECT 73.560 142.150 74.060 142.320 ;
        RECT 73.560 140.870 74.060 141.040 ;
        RECT 74.230 139.965 74.560 141.935 ;
        RECT 76.300 141.750 76.800 141.920 ;
        RECT 73.560 139.590 74.060 139.760 ;
        RECT 73.060 137.730 73.390 139.340 ;
        RECT 74.230 137.730 74.560 139.340 ;
        RECT 75.800 138.845 76.130 141.535 ;
        RECT 76.970 138.845 77.300 141.535 ;
        RECT 76.300 138.470 76.800 138.640 ;
        RECT 73.560 137.310 74.060 137.480 ;
        RECT 73.060 135.450 73.390 137.060 ;
        RECT 74.230 135.450 74.560 137.060 ;
        RECT 75.800 135.565 76.130 138.255 ;
        RECT 76.970 135.565 77.300 138.255 ;
        RECT 73.560 135.030 74.060 135.200 ;
        RECT 76.300 135.190 76.800 135.360 ;
        RECT 73.060 133.170 73.390 134.780 ;
        RECT 74.230 133.170 74.560 134.780 ;
        RECT 73.560 132.750 74.060 132.920 ;
        RECT 73.060 130.890 73.390 132.500 ;
        RECT 74.230 130.890 74.560 132.500 ;
        RECT 73.560 130.470 74.060 130.640 ;
        RECT 73.060 128.285 73.390 130.255 ;
        RECT 73.560 129.190 74.060 129.360 ;
        RECT 74.230 128.285 74.560 130.255 ;
        RECT 76.970 128.310 77.300 134.960 ;
        RECT 73.560 127.910 74.060 128.080 ;
        RECT 76.300 127.910 76.800 128.080 ;
        RECT 73.060 125.725 73.390 127.695 ;
        RECT 73.560 126.630 74.060 126.800 ;
        RECT 74.230 125.725 74.560 127.695 ;
        RECT 73.560 125.350 74.060 125.520 ;
        RECT 73.060 123.490 73.390 125.100 ;
        RECT 74.230 123.490 74.560 125.100 ;
        RECT 73.560 123.070 74.060 123.240 ;
        RECT 73.060 121.210 73.390 122.820 ;
        RECT 74.230 121.210 74.560 122.820 ;
        RECT 76.970 121.030 77.300 127.680 ;
        RECT 73.560 120.790 74.060 120.960 ;
        RECT 76.300 120.630 76.800 120.800 ;
        RECT 73.060 118.930 73.390 120.540 ;
        RECT 74.230 118.930 74.560 120.540 ;
        RECT 73.560 118.510 74.060 118.680 ;
        RECT 73.060 116.650 73.390 118.260 ;
        RECT 74.230 116.650 74.560 118.260 ;
        RECT 75.800 117.725 76.130 120.415 ;
        RECT 76.970 117.725 77.300 120.415 ;
        RECT 76.300 117.350 76.800 117.520 ;
        RECT 73.560 116.230 74.060 116.400 ;
        RECT 73.560 114.950 74.060 115.120 ;
        RECT 74.230 114.045 74.560 116.015 ;
        RECT 75.800 114.445 76.130 117.135 ;
        RECT 76.970 114.445 77.300 117.135 ;
        RECT 76.300 114.070 76.800 114.240 ;
        RECT 73.560 113.670 74.060 113.840 ;
        RECT 77.600 113.210 77.770 142.780 ;
        RECT 72.590 113.040 77.770 113.210 ;
        RECT 81.020 142.780 86.200 142.950 ;
        RECT 81.020 113.210 81.190 142.780 ;
        RECT 84.730 142.150 85.230 142.320 ;
        RECT 81.990 141.750 82.490 141.920 ;
        RECT 81.490 138.845 81.820 141.535 ;
        RECT 82.660 138.845 82.990 141.535 ;
        RECT 84.230 139.965 84.560 141.935 ;
        RECT 84.730 140.870 85.230 141.040 ;
        RECT 84.730 139.590 85.230 139.760 ;
        RECT 81.990 138.470 82.490 138.640 ;
        RECT 81.490 135.565 81.820 138.255 ;
        RECT 82.660 135.565 82.990 138.255 ;
        RECT 84.230 137.730 84.560 139.340 ;
        RECT 85.400 137.730 85.730 139.340 ;
        RECT 84.730 137.310 85.230 137.480 ;
        RECT 84.230 135.450 84.560 137.060 ;
        RECT 85.400 135.450 85.730 137.060 ;
        RECT 81.990 135.190 82.490 135.360 ;
        RECT 84.730 135.030 85.230 135.200 ;
        RECT 81.490 128.310 81.820 134.960 ;
        RECT 84.230 133.170 84.560 134.780 ;
        RECT 85.400 133.170 85.730 134.780 ;
        RECT 84.730 132.750 85.230 132.920 ;
        RECT 84.230 130.890 84.560 132.500 ;
        RECT 85.400 130.890 85.730 132.500 ;
        RECT 84.730 130.470 85.230 130.640 ;
        RECT 84.230 128.285 84.560 130.255 ;
        RECT 84.730 129.190 85.230 129.360 ;
        RECT 85.400 128.285 85.730 130.255 ;
        RECT 81.990 127.910 82.490 128.080 ;
        RECT 84.730 127.910 85.230 128.080 ;
        RECT 81.490 121.030 81.820 127.680 ;
        RECT 84.230 125.725 84.560 127.695 ;
        RECT 84.730 126.630 85.230 126.800 ;
        RECT 85.400 125.725 85.730 127.695 ;
        RECT 84.730 125.350 85.230 125.520 ;
        RECT 84.230 123.490 84.560 125.100 ;
        RECT 85.400 123.490 85.730 125.100 ;
        RECT 84.730 123.070 85.230 123.240 ;
        RECT 84.230 121.210 84.560 122.820 ;
        RECT 85.400 121.210 85.730 122.820 ;
        RECT 81.990 120.630 82.490 120.800 ;
        RECT 84.730 120.790 85.230 120.960 ;
        RECT 81.490 117.725 81.820 120.415 ;
        RECT 82.660 117.725 82.990 120.415 ;
        RECT 84.230 118.930 84.560 120.540 ;
        RECT 85.400 118.930 85.730 120.540 ;
        RECT 84.730 118.510 85.230 118.680 ;
        RECT 81.990 117.350 82.490 117.520 ;
        RECT 81.490 114.445 81.820 117.135 ;
        RECT 82.660 114.445 82.990 117.135 ;
        RECT 84.230 116.650 84.560 118.260 ;
        RECT 85.400 116.650 85.730 118.260 ;
        RECT 84.730 116.230 85.230 116.400 ;
        RECT 81.990 114.070 82.490 114.240 ;
        RECT 84.230 114.045 84.560 116.015 ;
        RECT 84.730 114.950 85.230 115.120 ;
        RECT 84.730 113.670 85.230 113.840 ;
        RECT 86.030 113.210 86.200 142.780 ;
        RECT 91.915 142.650 92.085 151.500 ;
        RECT 92.885 150.830 93.385 151.000 ;
        RECT 92.385 149.690 92.715 150.580 ;
        RECT 92.885 150.050 93.385 150.220 ;
        RECT 92.885 149.270 93.385 149.440 ;
        RECT 93.555 147.410 93.885 149.020 ;
        RECT 92.885 146.990 93.385 147.160 ;
        RECT 93.555 145.130 93.885 146.740 ;
        RECT 92.885 144.710 93.385 144.880 ;
        RECT 92.385 143.570 92.715 144.460 ;
        RECT 92.885 143.930 93.385 144.100 ;
        RECT 92.885 143.150 93.385 143.320 ;
        RECT 94.185 142.650 94.355 151.500 ;
        RECT 91.915 142.480 94.355 142.650 ;
        RECT 96.080 151.500 102.610 151.670 ;
        RECT 87.660 138.290 90.600 138.460 ;
        RECT 87.660 117.760 87.830 138.290 ;
        RECT 88.630 137.620 89.630 137.790 ;
        RECT 88.130 135.435 88.460 137.405 ;
        RECT 88.630 136.340 89.630 136.510 ;
        RECT 89.800 135.435 90.130 137.405 ;
        RECT 88.630 135.060 89.630 135.230 ;
        RECT 88.130 133.200 88.460 134.810 ;
        RECT 89.800 133.200 90.130 134.810 ;
        RECT 88.630 132.780 89.630 132.950 ;
        RECT 88.130 130.920 88.460 132.530 ;
        RECT 89.800 130.920 90.130 132.530 ;
        RECT 88.630 130.500 89.630 130.670 ;
        RECT 88.130 128.315 88.460 130.285 ;
        RECT 88.630 129.220 89.630 129.390 ;
        RECT 89.800 128.315 90.130 130.285 ;
        RECT 88.630 127.940 89.630 128.110 ;
        RECT 88.130 125.755 88.460 127.725 ;
        RECT 88.630 126.660 89.630 126.830 ;
        RECT 89.800 125.755 90.130 127.725 ;
        RECT 88.630 125.380 89.630 125.550 ;
        RECT 88.130 123.520 88.460 125.130 ;
        RECT 88.630 123.100 89.630 123.270 ;
        RECT 88.130 121.240 88.460 122.850 ;
        RECT 88.630 120.820 89.630 120.990 ;
        RECT 88.130 118.635 88.460 120.605 ;
        RECT 88.630 119.540 89.630 119.710 ;
        RECT 89.800 118.635 90.130 120.605 ;
        RECT 88.630 118.260 89.630 118.430 ;
        RECT 90.430 117.760 90.600 138.290 ;
        RECT 87.660 117.590 90.600 117.760 ;
        RECT 91.915 138.290 94.355 138.460 ;
        RECT 91.915 117.760 92.085 138.290 ;
        RECT 92.885 137.620 93.385 137.790 ;
        RECT 92.385 135.435 92.715 137.405 ;
        RECT 92.885 136.340 93.385 136.510 ;
        RECT 93.555 135.435 93.885 137.405 ;
        RECT 92.885 135.060 93.385 135.230 ;
        RECT 92.385 133.200 92.715 134.810 ;
        RECT 93.555 133.200 93.885 134.810 ;
        RECT 92.885 132.780 93.385 132.950 ;
        RECT 92.385 130.920 92.715 132.530 ;
        RECT 93.555 130.920 93.885 132.530 ;
        RECT 92.885 130.500 93.385 130.670 ;
        RECT 92.385 128.315 92.715 130.285 ;
        RECT 92.885 129.220 93.385 129.390 ;
        RECT 93.555 128.315 93.885 130.285 ;
        RECT 92.885 127.940 93.385 128.110 ;
        RECT 92.385 125.755 92.715 127.725 ;
        RECT 92.885 126.660 93.385 126.830 ;
        RECT 93.555 125.755 93.885 127.725 ;
        RECT 92.885 125.380 93.385 125.550 ;
        RECT 93.555 123.520 93.885 125.130 ;
        RECT 92.885 123.100 93.385 123.270 ;
        RECT 93.555 121.240 93.885 122.850 ;
        RECT 92.885 120.820 93.385 120.990 ;
        RECT 92.385 118.635 92.715 120.605 ;
        RECT 92.885 119.540 93.385 119.710 ;
        RECT 93.555 118.635 93.885 120.605 ;
        RECT 92.885 118.260 93.385 118.430 ;
        RECT 94.185 117.760 94.355 138.290 ;
        RECT 91.915 117.590 94.355 117.760 ;
        RECT 81.020 113.040 86.200 113.210 ;
        RECT 88.545 113.340 91.120 113.510 ;
        RECT 91.505 113.340 95.105 113.510 ;
        RECT 63.685 89.200 67.285 89.370 ;
        RECT 67.670 89.200 70.245 89.370 ;
        RECT 88.545 89.370 88.715 113.340 ;
        RECT 89.175 112.670 89.675 112.840 ;
        RECT 93.475 112.670 94.475 112.840 ;
        RECT 89.845 110.810 90.175 112.420 ;
        RECT 92.975 110.810 93.305 112.420 ;
        RECT 89.175 110.390 89.675 110.560 ;
        RECT 93.475 110.390 94.475 110.560 ;
        RECT 89.845 108.530 90.175 110.140 ;
        RECT 92.975 108.530 93.305 110.140 ;
        RECT 89.175 108.110 89.675 108.280 ;
        RECT 93.475 108.110 94.475 108.280 ;
        RECT 89.845 106.250 90.175 107.860 ;
        RECT 92.975 106.250 93.305 107.860 ;
        RECT 89.175 105.830 89.675 106.000 ;
        RECT 93.475 105.830 94.475 106.000 ;
        RECT 89.845 103.970 90.175 105.580 ;
        RECT 92.975 103.970 93.305 105.580 ;
        RECT 89.175 103.550 89.675 103.720 ;
        RECT 93.475 103.550 94.475 103.720 ;
        RECT 89.845 101.690 90.175 103.300 ;
        RECT 92.975 101.690 93.305 103.300 ;
        RECT 89.175 101.270 89.675 101.440 ;
        RECT 93.475 101.270 94.475 101.440 ;
        RECT 89.845 99.410 90.175 101.020 ;
        RECT 92.975 99.410 93.305 101.020 ;
        RECT 89.175 98.990 89.675 99.160 ;
        RECT 93.475 98.990 94.475 99.160 ;
        RECT 89.845 97.130 90.175 98.740 ;
        RECT 92.975 97.130 93.305 98.740 ;
        RECT 89.175 96.710 89.675 96.880 ;
        RECT 93.475 96.710 94.475 96.880 ;
        RECT 89.845 94.850 90.175 96.460 ;
        RECT 92.975 94.850 93.305 96.460 ;
        RECT 89.175 94.430 89.675 94.600 ;
        RECT 93.475 94.430 94.475 94.600 ;
        RECT 89.845 92.570 90.175 94.180 ;
        RECT 92.975 92.570 93.305 94.180 ;
        RECT 89.175 92.150 89.675 92.320 ;
        RECT 93.475 92.150 94.475 92.320 ;
        RECT 89.845 90.290 90.175 91.900 ;
        RECT 92.975 90.290 93.305 91.900 ;
        RECT 89.175 89.870 89.675 90.040 ;
        RECT 93.475 89.870 94.475 90.040 ;
        RECT 94.935 89.370 95.105 113.340 ;
        RECT 96.080 112.170 96.250 151.500 ;
        RECT 97.050 150.830 98.050 151.000 ;
        RECT 97.050 150.050 98.050 150.220 ;
        RECT 98.220 149.690 98.550 150.580 ;
        RECT 97.050 149.270 98.050 149.440 ;
        RECT 96.550 147.410 96.880 149.020 ;
        RECT 97.050 146.990 98.050 147.160 ;
        RECT 96.550 145.130 96.880 146.740 ;
        RECT 97.050 144.710 98.050 144.880 ;
        RECT 97.050 143.930 98.050 144.100 ;
        RECT 98.220 143.570 98.550 144.460 ;
        RECT 97.050 143.150 98.050 143.320 ;
        RECT 97.050 142.370 98.050 142.540 ;
        RECT 98.220 142.010 98.550 142.900 ;
        RECT 97.050 141.590 98.050 141.760 ;
        RECT 100.640 141.590 101.640 141.760 ;
        RECT 96.550 139.730 96.880 141.340 ;
        RECT 98.220 139.730 98.550 141.340 ;
        RECT 100.140 139.730 100.470 141.340 ;
        RECT 97.050 139.310 98.050 139.480 ;
        RECT 100.640 139.310 101.640 139.480 ;
        RECT 96.550 137.450 96.880 139.060 ;
        RECT 98.220 137.450 98.550 139.060 ;
        RECT 100.140 137.450 100.470 139.060 ;
        RECT 97.050 137.030 98.050 137.200 ;
        RECT 100.640 137.030 101.640 137.200 ;
        RECT 96.550 135.170 96.880 136.780 ;
        RECT 98.220 135.170 98.550 136.780 ;
        RECT 100.140 135.170 100.470 136.780 ;
        RECT 97.050 134.750 98.050 134.920 ;
        RECT 100.640 134.750 101.640 134.920 ;
        RECT 96.550 132.890 96.880 134.500 ;
        RECT 98.220 132.890 98.550 134.500 ;
        RECT 100.140 132.890 100.470 134.500 ;
        RECT 97.050 132.470 98.050 132.640 ;
        RECT 100.640 132.470 101.640 132.640 ;
        RECT 96.550 130.610 96.880 132.220 ;
        RECT 98.220 130.610 98.550 132.220 ;
        RECT 100.140 130.610 100.470 132.220 ;
        RECT 97.050 130.190 98.050 130.360 ;
        RECT 100.640 130.190 101.640 130.360 ;
        RECT 96.550 128.330 96.880 129.940 ;
        RECT 98.220 128.330 98.550 129.940 ;
        RECT 101.810 128.330 102.140 129.940 ;
        RECT 97.050 127.910 98.050 128.080 ;
        RECT 100.640 127.910 101.640 128.080 ;
        RECT 96.550 126.050 96.880 127.660 ;
        RECT 98.220 126.050 98.550 127.660 ;
        RECT 101.810 126.050 102.140 127.660 ;
        RECT 97.050 125.630 98.050 125.800 ;
        RECT 100.640 125.630 101.640 125.800 ;
        RECT 96.550 123.770 96.880 125.380 ;
        RECT 98.220 123.770 98.550 125.380 ;
        RECT 100.140 123.770 100.470 125.380 ;
        RECT 97.050 123.350 98.050 123.520 ;
        RECT 100.640 123.350 101.640 123.520 ;
        RECT 96.550 121.490 96.880 123.100 ;
        RECT 98.220 121.490 98.550 123.100 ;
        RECT 100.140 121.490 100.470 123.100 ;
        RECT 97.050 121.070 98.050 121.240 ;
        RECT 100.640 121.070 101.640 121.240 ;
        RECT 96.550 119.210 96.880 120.820 ;
        RECT 98.220 119.210 98.550 120.820 ;
        RECT 100.140 119.210 100.470 120.820 ;
        RECT 97.050 118.790 98.050 118.960 ;
        RECT 100.640 118.790 101.640 118.960 ;
        RECT 96.550 116.930 96.880 118.540 ;
        RECT 98.220 116.930 98.550 118.540 ;
        RECT 100.140 116.930 100.470 118.540 ;
        RECT 97.050 116.510 98.050 116.680 ;
        RECT 100.640 116.510 101.640 116.680 ;
        RECT 96.550 114.650 96.880 116.260 ;
        RECT 98.220 114.650 98.550 116.260 ;
        RECT 100.140 114.650 100.470 116.260 ;
        RECT 97.050 114.230 98.050 114.400 ;
        RECT 100.640 114.230 101.640 114.400 ;
        RECT 97.050 113.450 98.050 113.620 ;
        RECT 98.220 113.090 98.550 113.980 ;
        RECT 97.050 112.670 98.050 112.840 ;
        RECT 102.440 112.170 102.610 151.500 ;
        RECT 96.080 112.000 102.610 112.170 ;
        RECT 88.545 89.200 91.120 89.370 ;
        RECT 91.505 89.200 95.105 89.370 ;
        RECT 88.505 83.020 91.080 83.190 ;
        RECT 91.490 83.020 95.090 83.190 ;
        RECT 71.475 82.670 74.330 82.840 ;
        RECT 74.860 82.670 83.700 82.840 ;
        RECT 84.230 82.670 87.085 82.840 ;
        RECT 71.475 78.060 71.645 82.670 ;
        RECT 72.445 82.000 73.445 82.170 ;
        RECT 75.745 82.000 76.745 82.170 ;
        RECT 77.395 82.000 78.395 82.170 ;
        RECT 71.945 81.390 72.275 81.920 ;
        RECT 72.445 81.570 73.445 81.740 ;
        RECT 73.615 81.390 73.945 81.920 ;
        RECT 75.245 81.390 75.575 81.920 ;
        RECT 75.745 81.570 76.745 81.740 ;
        RECT 77.395 81.570 78.395 81.740 ;
        RECT 78.565 81.390 78.895 81.920 ;
        RECT 72.445 81.140 73.445 81.310 ;
        RECT 75.745 81.140 76.745 81.310 ;
        RECT 77.395 81.140 78.395 81.310 ;
        RECT 71.945 80.530 72.275 81.060 ;
        RECT 72.445 80.710 73.445 80.880 ;
        RECT 73.615 80.530 73.945 81.060 ;
        RECT 75.245 80.530 75.575 81.060 ;
        RECT 75.745 80.710 76.745 80.880 ;
        RECT 77.395 80.710 78.395 80.880 ;
        RECT 78.565 80.530 78.895 81.060 ;
        RECT 72.445 80.280 73.445 80.450 ;
        RECT 75.745 80.280 76.745 80.450 ;
        RECT 77.395 80.280 78.395 80.450 ;
        RECT 71.945 79.670 72.275 80.200 ;
        RECT 72.445 79.850 73.445 80.020 ;
        RECT 73.615 79.670 73.945 80.200 ;
        RECT 75.245 79.670 75.575 80.200 ;
        RECT 75.745 79.850 76.745 80.020 ;
        RECT 77.395 79.850 78.395 80.020 ;
        RECT 78.565 79.670 78.895 80.200 ;
        RECT 72.445 79.420 73.445 79.590 ;
        RECT 75.745 79.420 76.745 79.590 ;
        RECT 77.395 79.420 78.395 79.590 ;
        RECT 71.945 78.810 72.275 79.340 ;
        RECT 72.445 78.990 73.445 79.160 ;
        RECT 73.615 78.810 73.945 79.340 ;
        RECT 75.245 78.810 75.575 79.340 ;
        RECT 75.745 78.990 76.745 79.160 ;
        RECT 77.395 78.990 78.395 79.160 ;
        RECT 78.565 78.810 78.895 79.340 ;
        RECT 72.445 78.560 73.445 78.730 ;
        RECT 75.745 78.560 76.745 78.730 ;
        RECT 77.395 78.560 78.395 78.730 ;
        RECT 79.195 78.060 79.365 82.670 ;
        RECT 80.165 82.000 81.165 82.170 ;
        RECT 81.815 82.000 82.815 82.170 ;
        RECT 85.115 82.000 86.115 82.170 ;
        RECT 79.665 81.390 79.995 81.920 ;
        RECT 80.165 81.570 81.165 81.740 ;
        RECT 81.815 81.570 82.815 81.740 ;
        RECT 82.985 81.390 83.315 81.920 ;
        RECT 84.615 81.390 84.945 81.920 ;
        RECT 85.115 81.570 86.115 81.740 ;
        RECT 86.285 81.390 86.615 81.920 ;
        RECT 80.165 81.140 81.165 81.310 ;
        RECT 81.815 81.140 82.815 81.310 ;
        RECT 85.115 81.140 86.115 81.310 ;
        RECT 79.665 80.530 79.995 81.060 ;
        RECT 80.165 80.710 81.165 80.880 ;
        RECT 81.815 80.710 82.815 80.880 ;
        RECT 82.985 80.530 83.315 81.060 ;
        RECT 84.615 80.530 84.945 81.060 ;
        RECT 85.115 80.710 86.115 80.880 ;
        RECT 86.285 80.530 86.615 81.060 ;
        RECT 80.165 80.280 81.165 80.450 ;
        RECT 81.815 80.280 82.815 80.450 ;
        RECT 85.115 80.280 86.115 80.450 ;
        RECT 79.665 79.670 79.995 80.200 ;
        RECT 80.165 79.850 81.165 80.020 ;
        RECT 81.815 79.850 82.815 80.020 ;
        RECT 82.985 79.670 83.315 80.200 ;
        RECT 84.615 79.670 84.945 80.200 ;
        RECT 85.115 79.850 86.115 80.020 ;
        RECT 86.285 79.670 86.615 80.200 ;
        RECT 80.165 79.420 81.165 79.590 ;
        RECT 81.815 79.420 82.815 79.590 ;
        RECT 85.115 79.420 86.115 79.590 ;
        RECT 79.665 78.810 79.995 79.340 ;
        RECT 80.165 78.990 81.165 79.160 ;
        RECT 81.815 78.990 82.815 79.160 ;
        RECT 82.985 78.810 83.315 79.340 ;
        RECT 84.615 78.810 84.945 79.340 ;
        RECT 85.115 78.990 86.115 79.160 ;
        RECT 86.285 78.810 86.615 79.340 ;
        RECT 80.165 78.560 81.165 78.730 ;
        RECT 81.815 78.560 82.815 78.730 ;
        RECT 85.115 78.560 86.115 78.730 ;
        RECT 86.915 78.060 87.085 82.670 ;
        RECT 88.505 78.410 88.675 83.020 ;
        RECT 89.110 82.350 90.110 82.520 ;
        RECT 92.460 82.350 94.460 82.520 ;
        RECT 89.110 81.920 90.110 82.090 ;
        RECT 90.280 81.740 90.610 82.270 ;
        RECT 91.960 81.740 92.290 82.270 ;
        RECT 92.460 81.920 94.460 82.090 ;
        RECT 89.110 81.490 90.110 81.660 ;
        RECT 92.460 81.490 94.460 81.660 ;
        RECT 89.110 81.060 90.110 81.230 ;
        RECT 90.280 80.880 90.610 81.410 ;
        RECT 91.960 80.880 92.290 81.410 ;
        RECT 92.460 81.060 94.460 81.230 ;
        RECT 89.110 80.630 90.110 80.800 ;
        RECT 92.460 80.630 94.460 80.800 ;
        RECT 89.110 80.200 90.110 80.370 ;
        RECT 90.280 80.020 90.610 80.550 ;
        RECT 91.960 80.020 92.290 80.550 ;
        RECT 92.460 80.200 94.460 80.370 ;
        RECT 89.110 79.770 90.110 79.940 ;
        RECT 92.460 79.770 94.460 79.940 ;
        RECT 89.110 79.340 90.110 79.510 ;
        RECT 90.280 79.160 90.610 79.690 ;
        RECT 91.960 79.160 92.290 79.690 ;
        RECT 92.460 79.340 94.460 79.510 ;
        RECT 89.110 78.910 90.110 79.080 ;
        RECT 92.460 78.910 94.460 79.080 ;
        RECT 94.920 78.410 95.090 83.020 ;
        RECT 88.505 78.240 91.080 78.410 ;
        RECT 91.490 78.240 95.090 78.410 ;
        RECT 71.475 77.890 74.330 78.060 ;
        RECT 74.860 77.890 83.700 78.060 ;
        RECT 84.230 77.890 87.085 78.060 ;
        RECT 64.725 72.360 67.300 72.530 ;
        RECT 67.710 72.360 71.310 72.530 ;
        RECT 64.725 63.450 64.895 72.360 ;
        RECT 65.330 71.690 66.330 71.860 ;
        RECT 68.680 71.690 70.680 71.860 ;
        RECT 65.330 71.260 66.330 71.430 ;
        RECT 66.500 71.080 66.830 71.610 ;
        RECT 68.180 71.080 68.510 71.610 ;
        RECT 68.680 71.260 70.680 71.430 ;
        RECT 65.330 70.830 66.330 71.000 ;
        RECT 68.680 70.830 70.680 71.000 ;
        RECT 65.330 70.400 66.330 70.570 ;
        RECT 66.500 70.220 66.830 70.750 ;
        RECT 68.180 70.220 68.510 70.750 ;
        RECT 68.680 70.400 70.680 70.570 ;
        RECT 65.330 69.970 66.330 70.140 ;
        RECT 68.680 69.970 70.680 70.140 ;
        RECT 65.330 69.540 66.330 69.710 ;
        RECT 66.500 69.360 66.830 69.890 ;
        RECT 68.180 69.360 68.510 69.890 ;
        RECT 68.680 69.540 70.680 69.710 ;
        RECT 65.330 69.110 66.330 69.280 ;
        RECT 68.680 69.110 70.680 69.280 ;
        RECT 65.330 68.680 66.330 68.850 ;
        RECT 66.500 68.500 66.830 69.030 ;
        RECT 68.180 68.500 68.510 69.030 ;
        RECT 68.680 68.680 70.680 68.850 ;
        RECT 65.330 68.250 66.330 68.420 ;
        RECT 68.680 68.250 70.680 68.420 ;
        RECT 65.330 67.820 66.330 67.990 ;
        RECT 66.500 67.640 66.830 68.170 ;
        RECT 68.180 67.640 68.510 68.170 ;
        RECT 68.680 67.820 70.680 67.990 ;
        RECT 65.330 67.390 66.330 67.560 ;
        RECT 68.680 67.390 70.680 67.560 ;
        RECT 65.330 66.960 66.330 67.130 ;
        RECT 66.500 66.780 66.830 67.310 ;
        RECT 68.180 66.780 68.510 67.310 ;
        RECT 68.680 66.960 70.680 67.130 ;
        RECT 65.330 66.530 66.330 66.700 ;
        RECT 68.680 66.530 70.680 66.700 ;
        RECT 65.330 66.100 66.330 66.270 ;
        RECT 66.500 65.920 66.830 66.450 ;
        RECT 68.180 65.920 68.510 66.450 ;
        RECT 68.680 66.100 70.680 66.270 ;
        RECT 65.330 65.670 66.330 65.840 ;
        RECT 68.680 65.670 70.680 65.840 ;
        RECT 65.330 65.240 66.330 65.410 ;
        RECT 66.500 65.060 66.830 65.590 ;
        RECT 68.180 65.060 68.510 65.590 ;
        RECT 68.680 65.240 70.680 65.410 ;
        RECT 65.330 64.810 66.330 64.980 ;
        RECT 68.680 64.810 70.680 64.980 ;
        RECT 65.330 64.380 66.330 64.550 ;
        RECT 66.500 64.200 66.830 64.730 ;
        RECT 68.180 64.200 68.510 64.730 ;
        RECT 68.680 64.380 70.680 64.550 ;
        RECT 65.330 63.950 66.330 64.120 ;
        RECT 68.680 63.950 70.680 64.120 ;
        RECT 71.140 63.450 71.310 72.360 ;
        RECT 64.725 63.280 67.300 63.450 ;
        RECT 67.710 63.280 71.310 63.450 ;
        RECT 73.745 72.360 76.320 72.530 ;
        RECT 76.730 72.360 83.760 72.530 ;
        RECT 84.170 72.360 86.745 72.530 ;
        RECT 73.745 63.450 73.915 72.360 ;
        RECT 74.350 71.690 75.350 71.860 ;
        RECT 77.700 71.690 79.700 71.860 ;
        RECT 74.350 71.260 75.350 71.430 ;
        RECT 75.520 71.080 75.850 71.610 ;
        RECT 77.200 71.080 77.530 71.610 ;
        RECT 77.700 71.260 79.700 71.430 ;
        RECT 74.350 70.830 75.350 71.000 ;
        RECT 77.700 70.830 79.700 71.000 ;
        RECT 74.350 70.400 75.350 70.570 ;
        RECT 75.520 70.220 75.850 70.750 ;
        RECT 77.200 70.220 77.530 70.750 ;
        RECT 77.700 70.400 79.700 70.570 ;
        RECT 74.350 69.970 75.350 70.140 ;
        RECT 77.700 69.970 79.700 70.140 ;
        RECT 74.350 69.540 75.350 69.710 ;
        RECT 75.520 69.360 75.850 69.890 ;
        RECT 77.200 69.360 77.530 69.890 ;
        RECT 77.700 69.540 79.700 69.710 ;
        RECT 74.350 69.110 75.350 69.280 ;
        RECT 77.700 69.110 79.700 69.280 ;
        RECT 74.350 68.680 75.350 68.850 ;
        RECT 75.520 68.500 75.850 69.030 ;
        RECT 77.200 68.500 77.530 69.030 ;
        RECT 77.700 68.680 79.700 68.850 ;
        RECT 74.350 68.250 75.350 68.420 ;
        RECT 77.700 68.250 79.700 68.420 ;
        RECT 74.350 67.820 75.350 67.990 ;
        RECT 75.520 67.640 75.850 68.170 ;
        RECT 77.200 67.640 77.530 68.170 ;
        RECT 77.700 67.820 79.700 67.990 ;
        RECT 74.350 67.390 75.350 67.560 ;
        RECT 77.700 67.390 79.700 67.560 ;
        RECT 74.350 66.960 75.350 67.130 ;
        RECT 75.520 66.780 75.850 67.310 ;
        RECT 77.200 66.780 77.530 67.310 ;
        RECT 77.700 66.960 79.700 67.130 ;
        RECT 74.350 66.530 75.350 66.700 ;
        RECT 77.700 66.530 79.700 66.700 ;
        RECT 74.350 66.100 75.350 66.270 ;
        RECT 75.520 65.920 75.850 66.450 ;
        RECT 77.200 65.920 77.530 66.450 ;
        RECT 77.700 66.100 79.700 66.270 ;
        RECT 74.350 65.670 75.350 65.840 ;
        RECT 77.700 65.670 79.700 65.840 ;
        RECT 74.350 65.240 75.350 65.410 ;
        RECT 75.520 65.060 75.850 65.590 ;
        RECT 77.200 65.060 77.530 65.590 ;
        RECT 77.700 65.240 79.700 65.410 ;
        RECT 74.350 64.810 75.350 64.980 ;
        RECT 77.700 64.810 79.700 64.980 ;
        RECT 74.350 64.380 75.350 64.550 ;
        RECT 75.520 64.200 75.850 64.730 ;
        RECT 77.200 64.200 77.530 64.730 ;
        RECT 77.700 64.380 79.700 64.550 ;
        RECT 74.350 63.950 75.350 64.120 ;
        RECT 77.700 63.950 79.700 64.120 ;
        RECT 80.160 63.450 80.330 72.360 ;
        RECT 80.790 71.690 82.790 71.860 ;
        RECT 85.140 71.690 86.140 71.860 ;
        RECT 80.790 71.260 82.790 71.430 ;
        RECT 82.960 71.080 83.290 71.610 ;
        RECT 84.640 71.080 84.970 71.610 ;
        RECT 85.140 71.260 86.140 71.430 ;
        RECT 80.790 70.830 82.790 71.000 ;
        RECT 85.140 70.830 86.140 71.000 ;
        RECT 80.790 70.400 82.790 70.570 ;
        RECT 82.960 70.220 83.290 70.750 ;
        RECT 84.640 70.220 84.970 70.750 ;
        RECT 85.140 70.400 86.140 70.570 ;
        RECT 80.790 69.970 82.790 70.140 ;
        RECT 85.140 69.970 86.140 70.140 ;
        RECT 80.790 69.540 82.790 69.710 ;
        RECT 82.960 69.360 83.290 69.890 ;
        RECT 84.640 69.360 84.970 69.890 ;
        RECT 85.140 69.540 86.140 69.710 ;
        RECT 80.790 69.110 82.790 69.280 ;
        RECT 85.140 69.110 86.140 69.280 ;
        RECT 80.790 68.680 82.790 68.850 ;
        RECT 82.960 68.500 83.290 69.030 ;
        RECT 84.640 68.500 84.970 69.030 ;
        RECT 85.140 68.680 86.140 68.850 ;
        RECT 80.790 68.250 82.790 68.420 ;
        RECT 85.140 68.250 86.140 68.420 ;
        RECT 80.790 67.820 82.790 67.990 ;
        RECT 82.960 67.640 83.290 68.170 ;
        RECT 84.640 67.640 84.970 68.170 ;
        RECT 85.140 67.820 86.140 67.990 ;
        RECT 80.790 67.390 82.790 67.560 ;
        RECT 85.140 67.390 86.140 67.560 ;
        RECT 80.790 66.960 82.790 67.130 ;
        RECT 82.960 66.780 83.290 67.310 ;
        RECT 84.640 66.780 84.970 67.310 ;
        RECT 85.140 66.960 86.140 67.130 ;
        RECT 80.790 66.530 82.790 66.700 ;
        RECT 85.140 66.530 86.140 66.700 ;
        RECT 80.790 66.100 82.790 66.270 ;
        RECT 82.960 65.920 83.290 66.450 ;
        RECT 84.640 65.920 84.970 66.450 ;
        RECT 85.140 66.100 86.140 66.270 ;
        RECT 80.790 65.670 82.790 65.840 ;
        RECT 85.140 65.670 86.140 65.840 ;
        RECT 80.790 65.240 82.790 65.410 ;
        RECT 82.960 65.060 83.290 65.590 ;
        RECT 84.640 65.060 84.970 65.590 ;
        RECT 85.140 65.240 86.140 65.410 ;
        RECT 80.790 64.810 82.790 64.980 ;
        RECT 85.140 64.810 86.140 64.980 ;
        RECT 80.790 64.380 82.790 64.550 ;
        RECT 82.960 64.200 83.290 64.730 ;
        RECT 84.640 64.200 84.970 64.730 ;
        RECT 85.140 64.380 86.140 64.550 ;
        RECT 80.790 63.950 82.790 64.120 ;
        RECT 85.140 63.950 86.140 64.120 ;
        RECT 86.575 63.450 86.745 72.360 ;
        RECT 73.745 63.280 76.320 63.450 ;
        RECT 76.730 63.280 83.760 63.450 ;
        RECT 84.170 63.280 86.745 63.450 ;
        RECT 88.505 72.360 91.080 72.530 ;
        RECT 91.490 72.360 95.090 72.530 ;
        RECT 88.505 63.450 88.675 72.360 ;
        RECT 89.110 71.690 90.110 71.860 ;
        RECT 92.460 71.690 94.460 71.860 ;
        RECT 89.110 71.260 90.110 71.430 ;
        RECT 90.280 71.080 90.610 71.610 ;
        RECT 91.960 71.080 92.290 71.610 ;
        RECT 92.460 71.260 94.460 71.430 ;
        RECT 89.110 70.830 90.110 71.000 ;
        RECT 92.460 70.830 94.460 71.000 ;
        RECT 89.110 70.400 90.110 70.570 ;
        RECT 90.280 70.220 90.610 70.750 ;
        RECT 91.960 70.220 92.290 70.750 ;
        RECT 92.460 70.400 94.460 70.570 ;
        RECT 89.110 69.970 90.110 70.140 ;
        RECT 92.460 69.970 94.460 70.140 ;
        RECT 89.110 69.540 90.110 69.710 ;
        RECT 90.280 69.360 90.610 69.890 ;
        RECT 91.960 69.360 92.290 69.890 ;
        RECT 92.460 69.540 94.460 69.710 ;
        RECT 89.110 69.110 90.110 69.280 ;
        RECT 92.460 69.110 94.460 69.280 ;
        RECT 89.110 68.680 90.110 68.850 ;
        RECT 90.280 68.500 90.610 69.030 ;
        RECT 91.960 68.500 92.290 69.030 ;
        RECT 92.460 68.680 94.460 68.850 ;
        RECT 89.110 68.250 90.110 68.420 ;
        RECT 92.460 68.250 94.460 68.420 ;
        RECT 89.110 67.820 90.110 67.990 ;
        RECT 90.280 67.640 90.610 68.170 ;
        RECT 91.960 67.640 92.290 68.170 ;
        RECT 92.460 67.820 94.460 67.990 ;
        RECT 89.110 67.390 90.110 67.560 ;
        RECT 92.460 67.390 94.460 67.560 ;
        RECT 89.110 66.960 90.110 67.130 ;
        RECT 90.280 66.780 90.610 67.310 ;
        RECT 91.960 66.780 92.290 67.310 ;
        RECT 92.460 66.960 94.460 67.130 ;
        RECT 89.110 66.530 90.110 66.700 ;
        RECT 92.460 66.530 94.460 66.700 ;
        RECT 89.110 66.100 90.110 66.270 ;
        RECT 90.280 65.920 90.610 66.450 ;
        RECT 91.960 65.920 92.290 66.450 ;
        RECT 92.460 66.100 94.460 66.270 ;
        RECT 89.110 65.670 90.110 65.840 ;
        RECT 92.460 65.670 94.460 65.840 ;
        RECT 89.110 65.240 90.110 65.410 ;
        RECT 90.280 65.060 90.610 65.590 ;
        RECT 91.960 65.060 92.290 65.590 ;
        RECT 92.460 65.240 94.460 65.410 ;
        RECT 89.110 64.810 90.110 64.980 ;
        RECT 92.460 64.810 94.460 64.980 ;
        RECT 89.110 64.380 90.110 64.550 ;
        RECT 90.280 64.200 90.610 64.730 ;
        RECT 91.960 64.200 92.290 64.730 ;
        RECT 92.460 64.380 94.460 64.550 ;
        RECT 89.110 63.950 90.110 64.120 ;
        RECT 92.460 63.950 94.460 64.120 ;
        RECT 94.920 63.450 95.090 72.360 ;
        RECT 88.505 63.280 91.080 63.450 ;
        RECT 91.490 63.280 95.090 63.450 ;
        RECT 108.635 63.260 108.805 164.750 ;
        RECT 109.605 164.080 110.305 164.250 ;
        RECT 110.975 164.080 111.675 164.250 ;
        RECT 112.345 164.080 113.045 164.250 ;
        RECT 110.475 162.220 110.805 163.830 ;
        RECT 111.845 162.220 112.175 163.830 ;
        RECT 109.605 161.800 110.305 161.970 ;
        RECT 110.975 161.800 111.675 161.970 ;
        RECT 112.345 161.800 113.045 161.970 ;
        RECT 110.475 159.940 110.805 161.550 ;
        RECT 111.845 159.940 112.175 161.550 ;
        RECT 109.605 159.520 110.305 159.690 ;
        RECT 110.975 159.520 111.675 159.690 ;
        RECT 112.345 159.520 113.045 159.690 ;
        RECT 110.475 157.660 110.805 159.270 ;
        RECT 111.845 157.660 112.175 159.270 ;
        RECT 109.605 157.240 110.305 157.410 ;
        RECT 110.975 157.240 111.675 157.410 ;
        RECT 112.345 157.240 113.045 157.410 ;
        RECT 110.475 155.380 110.805 156.990 ;
        RECT 111.845 155.380 112.175 156.990 ;
        RECT 109.605 154.960 110.305 155.130 ;
        RECT 110.975 154.960 111.675 155.130 ;
        RECT 112.345 154.960 113.045 155.130 ;
        RECT 110.475 153.100 110.805 154.710 ;
        RECT 111.845 153.100 112.175 154.710 ;
        RECT 109.605 152.680 110.305 152.850 ;
        RECT 110.975 152.680 111.675 152.850 ;
        RECT 112.345 152.680 113.045 152.850 ;
        RECT 110.475 150.820 110.805 152.430 ;
        RECT 111.845 150.820 112.175 152.430 ;
        RECT 109.605 150.400 110.305 150.570 ;
        RECT 110.975 150.400 111.675 150.570 ;
        RECT 112.345 150.400 113.045 150.570 ;
        RECT 110.475 148.540 110.805 150.150 ;
        RECT 111.845 148.540 112.175 150.150 ;
        RECT 109.605 148.120 110.305 148.290 ;
        RECT 110.975 148.120 111.675 148.290 ;
        RECT 112.345 148.120 113.045 148.290 ;
        RECT 110.475 146.260 110.805 147.870 ;
        RECT 111.845 146.260 112.175 147.870 ;
        RECT 109.605 145.840 110.305 146.010 ;
        RECT 110.975 145.840 111.675 146.010 ;
        RECT 112.345 145.840 113.045 146.010 ;
        RECT 110.475 143.980 110.805 145.590 ;
        RECT 111.845 143.980 112.175 145.590 ;
        RECT 109.605 143.560 110.305 143.730 ;
        RECT 110.975 143.560 111.675 143.730 ;
        RECT 112.345 143.560 113.045 143.730 ;
        RECT 110.475 141.700 110.805 143.310 ;
        RECT 111.845 141.700 112.175 143.310 ;
        RECT 109.605 141.280 110.305 141.450 ;
        RECT 110.975 141.280 111.675 141.450 ;
        RECT 112.345 141.280 113.045 141.450 ;
        RECT 110.475 139.420 110.805 141.030 ;
        RECT 111.845 139.420 112.175 141.030 ;
        RECT 109.605 139.000 110.305 139.170 ;
        RECT 110.975 139.000 111.675 139.170 ;
        RECT 112.345 139.000 113.045 139.170 ;
        RECT 110.475 137.140 110.805 138.750 ;
        RECT 111.845 137.140 112.175 138.750 ;
        RECT 109.605 136.720 110.305 136.890 ;
        RECT 110.975 136.720 111.675 136.890 ;
        RECT 112.345 136.720 113.045 136.890 ;
        RECT 110.475 134.860 110.805 136.470 ;
        RECT 111.845 134.860 112.175 136.470 ;
        RECT 109.605 134.440 110.305 134.610 ;
        RECT 110.975 134.440 111.675 134.610 ;
        RECT 112.345 134.440 113.045 134.610 ;
        RECT 110.475 132.580 110.805 134.190 ;
        RECT 111.845 132.580 112.175 134.190 ;
        RECT 109.605 132.160 110.305 132.330 ;
        RECT 110.975 132.160 111.675 132.330 ;
        RECT 112.345 132.160 113.045 132.330 ;
        RECT 110.475 130.300 110.805 131.910 ;
        RECT 111.845 130.300 112.175 131.910 ;
        RECT 109.605 129.880 110.305 130.050 ;
        RECT 110.975 129.880 111.675 130.050 ;
        RECT 112.345 129.880 113.045 130.050 ;
        RECT 110.475 128.020 110.805 129.630 ;
        RECT 111.845 128.020 112.175 129.630 ;
        RECT 109.605 127.600 110.305 127.770 ;
        RECT 110.975 127.600 111.675 127.770 ;
        RECT 112.345 127.600 113.045 127.770 ;
        RECT 110.475 125.740 110.805 127.350 ;
        RECT 111.845 125.740 112.175 127.350 ;
        RECT 109.605 125.320 110.305 125.490 ;
        RECT 110.975 125.320 111.675 125.490 ;
        RECT 112.345 125.320 113.045 125.490 ;
        RECT 110.475 123.460 110.805 125.070 ;
        RECT 111.845 123.460 112.175 125.070 ;
        RECT 109.605 123.040 110.305 123.210 ;
        RECT 110.975 123.040 111.675 123.210 ;
        RECT 112.345 123.040 113.045 123.210 ;
        RECT 110.475 121.180 110.805 122.790 ;
        RECT 111.845 121.180 112.175 122.790 ;
        RECT 109.605 120.760 110.305 120.930 ;
        RECT 110.975 120.760 111.675 120.930 ;
        RECT 112.345 120.760 113.045 120.930 ;
        RECT 110.475 118.900 110.805 120.510 ;
        RECT 111.845 118.900 112.175 120.510 ;
        RECT 109.605 118.480 110.305 118.650 ;
        RECT 110.975 118.480 111.675 118.650 ;
        RECT 112.345 118.480 113.045 118.650 ;
        RECT 110.475 116.620 110.805 118.230 ;
        RECT 111.845 116.620 112.175 118.230 ;
        RECT 109.605 116.200 110.305 116.370 ;
        RECT 110.975 116.200 111.675 116.370 ;
        RECT 112.345 116.200 113.045 116.370 ;
        RECT 110.475 114.340 110.805 115.950 ;
        RECT 111.845 114.340 112.175 115.950 ;
        RECT 109.605 113.920 110.305 114.090 ;
        RECT 110.975 113.920 111.675 114.090 ;
        RECT 112.345 113.920 113.045 114.090 ;
        RECT 110.475 112.060 110.805 113.670 ;
        RECT 111.845 112.060 112.175 113.670 ;
        RECT 109.605 111.640 110.305 111.810 ;
        RECT 110.975 111.640 111.675 111.810 ;
        RECT 112.345 111.640 113.045 111.810 ;
        RECT 110.475 109.780 110.805 111.390 ;
        RECT 111.845 109.780 112.175 111.390 ;
        RECT 109.605 109.360 110.305 109.530 ;
        RECT 110.975 109.360 111.675 109.530 ;
        RECT 112.345 109.360 113.045 109.530 ;
        RECT 110.475 107.500 110.805 109.110 ;
        RECT 111.845 107.500 112.175 109.110 ;
        RECT 109.605 107.080 110.305 107.250 ;
        RECT 110.975 107.080 111.675 107.250 ;
        RECT 112.345 107.080 113.045 107.250 ;
        RECT 110.475 105.220 110.805 106.830 ;
        RECT 111.845 105.220 112.175 106.830 ;
        RECT 109.605 104.800 110.305 104.970 ;
        RECT 110.975 104.800 111.675 104.970 ;
        RECT 112.345 104.800 113.045 104.970 ;
        RECT 110.475 102.940 110.805 104.550 ;
        RECT 111.845 102.940 112.175 104.550 ;
        RECT 109.605 102.520 110.305 102.690 ;
        RECT 110.975 102.520 111.675 102.690 ;
        RECT 112.345 102.520 113.045 102.690 ;
        RECT 110.475 100.660 110.805 102.270 ;
        RECT 111.845 100.660 112.175 102.270 ;
        RECT 109.605 100.240 110.305 100.410 ;
        RECT 110.975 100.240 111.675 100.410 ;
        RECT 112.345 100.240 113.045 100.410 ;
        RECT 110.475 98.380 110.805 99.990 ;
        RECT 111.845 98.380 112.175 99.990 ;
        RECT 109.605 97.960 110.305 98.130 ;
        RECT 110.975 97.960 111.675 98.130 ;
        RECT 112.345 97.960 113.045 98.130 ;
        RECT 110.475 96.100 110.805 97.710 ;
        RECT 111.845 96.100 112.175 97.710 ;
        RECT 109.605 95.680 110.305 95.850 ;
        RECT 110.975 95.680 111.675 95.850 ;
        RECT 112.345 95.680 113.045 95.850 ;
        RECT 110.475 93.820 110.805 95.430 ;
        RECT 111.845 93.820 112.175 95.430 ;
        RECT 109.605 93.400 110.305 93.570 ;
        RECT 110.975 93.400 111.675 93.570 ;
        RECT 112.345 93.400 113.045 93.570 ;
        RECT 110.475 91.540 110.805 93.150 ;
        RECT 111.845 91.540 112.175 93.150 ;
        RECT 109.605 91.120 110.305 91.290 ;
        RECT 110.975 91.120 111.675 91.290 ;
        RECT 112.345 91.120 113.045 91.290 ;
        RECT 110.475 89.260 110.805 90.870 ;
        RECT 111.845 89.260 112.175 90.870 ;
        RECT 109.605 88.840 110.305 89.010 ;
        RECT 110.975 88.840 111.675 89.010 ;
        RECT 112.345 88.840 113.045 89.010 ;
        RECT 110.475 86.980 110.805 88.590 ;
        RECT 111.845 86.980 112.175 88.590 ;
        RECT 109.605 86.560 110.305 86.730 ;
        RECT 110.975 86.560 111.675 86.730 ;
        RECT 112.345 86.560 113.045 86.730 ;
        RECT 110.475 84.700 110.805 86.310 ;
        RECT 111.845 84.700 112.175 86.310 ;
        RECT 109.605 84.280 110.305 84.450 ;
        RECT 110.975 84.280 111.675 84.450 ;
        RECT 112.345 84.280 113.045 84.450 ;
        RECT 110.475 82.420 110.805 84.030 ;
        RECT 111.845 82.420 112.175 84.030 ;
        RECT 109.605 82.000 110.305 82.170 ;
        RECT 110.975 82.000 111.675 82.170 ;
        RECT 112.345 82.000 113.045 82.170 ;
        RECT 110.475 80.140 110.805 81.750 ;
        RECT 111.845 80.140 112.175 81.750 ;
        RECT 109.605 79.720 110.305 79.890 ;
        RECT 110.975 79.720 111.675 79.890 ;
        RECT 112.345 79.720 113.045 79.890 ;
        RECT 110.475 77.860 110.805 79.470 ;
        RECT 111.845 77.860 112.175 79.470 ;
        RECT 109.605 77.440 110.305 77.610 ;
        RECT 110.975 77.440 111.675 77.610 ;
        RECT 112.345 77.440 113.045 77.610 ;
        RECT 110.475 75.580 110.805 77.190 ;
        RECT 111.845 75.580 112.175 77.190 ;
        RECT 109.605 75.160 110.305 75.330 ;
        RECT 110.975 75.160 111.675 75.330 ;
        RECT 112.345 75.160 113.045 75.330 ;
        RECT 110.475 73.300 110.805 74.910 ;
        RECT 111.845 73.300 112.175 74.910 ;
        RECT 109.605 72.880 110.305 73.050 ;
        RECT 110.975 72.880 111.675 73.050 ;
        RECT 112.345 72.880 113.045 73.050 ;
        RECT 110.475 71.020 110.805 72.630 ;
        RECT 111.845 71.020 112.175 72.630 ;
        RECT 109.605 70.600 110.305 70.770 ;
        RECT 110.975 70.600 111.675 70.770 ;
        RECT 112.345 70.600 113.045 70.770 ;
        RECT 110.475 68.740 110.805 70.350 ;
        RECT 111.845 68.740 112.175 70.350 ;
        RECT 109.605 68.320 110.305 68.490 ;
        RECT 110.975 68.320 111.675 68.490 ;
        RECT 112.345 68.320 113.045 68.490 ;
        RECT 110.475 66.460 110.805 68.070 ;
        RECT 111.845 66.460 112.175 68.070 ;
        RECT 109.605 66.040 110.305 66.210 ;
        RECT 110.975 66.040 111.675 66.210 ;
        RECT 112.345 66.040 113.045 66.210 ;
        RECT 110.475 64.180 110.805 65.790 ;
        RECT 111.845 64.180 112.175 65.790 ;
        RECT 109.605 63.760 110.305 63.930 ;
        RECT 110.975 63.760 111.675 63.930 ;
        RECT 112.345 63.760 113.045 63.930 ;
        RECT 113.845 63.260 114.015 164.750 ;
        RECT 121.840 164.710 125.850 164.880 ;
        RECT 114.925 118.155 117.565 118.325 ;
        RECT 114.925 114.485 115.095 118.155 ;
        RECT 115.895 117.525 116.595 117.695 ;
        RECT 115.895 117.095 116.595 117.265 ;
        RECT 116.765 117.095 117.095 117.265 ;
        RECT 115.895 116.665 116.595 116.835 ;
        RECT 115.395 116.235 115.725 116.405 ;
        RECT 115.895 116.235 116.595 116.405 ;
        RECT 115.895 115.805 116.595 115.975 ;
        RECT 115.895 115.375 116.595 115.545 ;
        RECT 116.765 115.375 117.095 115.545 ;
        RECT 115.895 114.945 116.595 115.115 ;
        RECT 117.395 114.485 117.565 118.155 ;
        RECT 114.925 114.315 117.565 114.485 ;
        RECT 118.195 117.920 121.135 118.090 ;
        RECT 114.925 113.525 117.565 113.695 ;
        RECT 114.925 109.775 115.095 113.525 ;
        RECT 115.895 112.855 116.595 113.025 ;
        RECT 115.395 112.425 115.725 112.595 ;
        RECT 115.895 112.425 116.595 112.595 ;
        RECT 115.895 111.995 116.595 112.165 ;
        RECT 115.895 111.565 116.595 111.735 ;
        RECT 116.765 111.565 117.095 111.735 ;
        RECT 115.895 111.135 116.595 111.305 ;
        RECT 115.395 110.705 115.725 110.875 ;
        RECT 115.895 110.705 116.595 110.875 ;
        RECT 115.895 110.275 116.595 110.445 ;
        RECT 117.395 109.775 117.565 113.525 ;
        RECT 118.195 109.950 118.365 117.920 ;
        RECT 119.165 117.290 120.165 117.460 ;
        RECT 118.665 116.860 118.995 117.030 ;
        RECT 119.165 116.860 120.165 117.030 ;
        RECT 119.165 116.430 120.165 116.600 ;
        RECT 118.665 116.000 118.995 116.170 ;
        RECT 119.165 116.000 120.165 116.170 ;
        RECT 119.165 115.570 120.165 115.740 ;
        RECT 118.665 115.140 118.995 115.310 ;
        RECT 119.165 115.140 120.165 115.310 ;
        RECT 119.165 114.710 120.165 114.880 ;
        RECT 119.165 114.280 120.165 114.450 ;
        RECT 120.335 114.280 120.665 114.450 ;
        RECT 119.165 113.850 120.165 114.020 ;
        RECT 119.165 113.420 120.165 113.590 ;
        RECT 120.335 113.420 120.665 113.590 ;
        RECT 119.165 112.990 120.165 113.160 ;
        RECT 118.665 112.560 118.995 112.730 ;
        RECT 119.165 112.560 120.165 112.730 ;
        RECT 119.165 112.130 120.165 112.300 ;
        RECT 118.665 111.700 118.995 111.870 ;
        RECT 119.165 111.700 120.165 111.870 ;
        RECT 119.165 111.270 120.165 111.440 ;
        RECT 118.665 110.840 118.995 111.010 ;
        RECT 119.165 110.840 120.165 111.010 ;
        RECT 119.165 110.410 120.165 110.580 ;
        RECT 120.965 109.950 121.135 117.920 ;
        RECT 118.195 109.780 121.135 109.950 ;
        RECT 114.925 109.605 117.565 109.775 ;
        RECT 114.925 83.955 117.565 84.125 ;
        RECT 114.925 80.285 115.095 83.955 ;
        RECT 115.895 83.325 116.595 83.495 ;
        RECT 115.895 82.895 116.595 83.065 ;
        RECT 116.765 82.895 117.095 83.065 ;
        RECT 115.895 82.465 116.595 82.635 ;
        RECT 115.395 82.035 115.725 82.205 ;
        RECT 115.895 82.035 116.595 82.205 ;
        RECT 115.895 81.605 116.595 81.775 ;
        RECT 115.895 81.175 116.595 81.345 ;
        RECT 116.765 81.175 117.095 81.345 ;
        RECT 115.895 80.745 116.595 80.915 ;
        RECT 117.395 80.285 117.565 83.955 ;
        RECT 114.925 80.115 117.565 80.285 ;
        RECT 118.195 83.720 121.135 83.890 ;
        RECT 114.925 79.325 117.565 79.495 ;
        RECT 114.925 75.575 115.095 79.325 ;
        RECT 115.895 78.655 116.595 78.825 ;
        RECT 115.395 78.225 115.725 78.395 ;
        RECT 115.895 78.225 116.595 78.395 ;
        RECT 115.895 77.795 116.595 77.965 ;
        RECT 115.895 77.365 116.595 77.535 ;
        RECT 116.765 77.365 117.095 77.535 ;
        RECT 115.895 76.935 116.595 77.105 ;
        RECT 115.395 76.505 115.725 76.675 ;
        RECT 115.895 76.505 116.595 76.675 ;
        RECT 115.895 76.075 116.595 76.245 ;
        RECT 117.395 75.575 117.565 79.325 ;
        RECT 118.195 75.750 118.365 83.720 ;
        RECT 119.165 83.090 120.165 83.260 ;
        RECT 118.665 82.660 118.995 82.830 ;
        RECT 119.165 82.660 120.165 82.830 ;
        RECT 119.165 82.230 120.165 82.400 ;
        RECT 118.665 81.800 118.995 81.970 ;
        RECT 119.165 81.800 120.165 81.970 ;
        RECT 119.165 81.370 120.165 81.540 ;
        RECT 118.665 80.940 118.995 81.110 ;
        RECT 119.165 80.940 120.165 81.110 ;
        RECT 119.165 80.510 120.165 80.680 ;
        RECT 119.165 80.080 120.165 80.250 ;
        RECT 120.335 80.080 120.665 80.250 ;
        RECT 119.165 79.650 120.165 79.820 ;
        RECT 119.165 79.220 120.165 79.390 ;
        RECT 120.335 79.220 120.665 79.390 ;
        RECT 119.165 78.790 120.165 78.960 ;
        RECT 118.665 78.360 118.995 78.530 ;
        RECT 119.165 78.360 120.165 78.530 ;
        RECT 119.165 77.930 120.165 78.100 ;
        RECT 118.665 77.500 118.995 77.670 ;
        RECT 119.165 77.500 120.165 77.670 ;
        RECT 119.165 77.070 120.165 77.240 ;
        RECT 118.665 76.640 118.995 76.810 ;
        RECT 119.165 76.640 120.165 76.810 ;
        RECT 119.165 76.210 120.165 76.380 ;
        RECT 120.965 75.750 121.135 83.720 ;
        RECT 121.840 76.980 122.010 164.710 ;
        RECT 122.810 164.080 123.510 164.250 ;
        RECT 124.180 164.080 124.880 164.250 ;
        RECT 122.310 162.220 122.640 163.830 ;
        RECT 125.050 162.220 125.380 163.830 ;
        RECT 122.810 161.800 123.510 161.970 ;
        RECT 124.180 161.800 124.880 161.970 ;
        RECT 122.310 159.940 122.640 161.550 ;
        RECT 125.050 159.940 125.380 161.550 ;
        RECT 122.810 159.520 123.510 159.690 ;
        RECT 124.180 159.520 124.880 159.690 ;
        RECT 122.310 157.660 122.640 159.270 ;
        RECT 123.680 157.660 124.010 159.270 ;
        RECT 125.050 157.660 125.380 159.270 ;
        RECT 122.810 157.240 123.510 157.410 ;
        RECT 124.180 157.240 124.880 157.410 ;
        RECT 122.310 155.380 122.640 156.990 ;
        RECT 123.680 155.380 124.010 156.990 ;
        RECT 125.050 155.380 125.380 156.990 ;
        RECT 122.810 154.960 123.510 155.130 ;
        RECT 124.180 154.960 124.880 155.130 ;
        RECT 122.310 153.100 122.640 154.710 ;
        RECT 123.680 153.100 124.010 154.710 ;
        RECT 125.050 153.100 125.380 154.710 ;
        RECT 122.810 152.680 123.510 152.850 ;
        RECT 124.180 152.680 124.880 152.850 ;
        RECT 122.310 150.820 122.640 152.430 ;
        RECT 123.680 150.820 124.010 152.430 ;
        RECT 125.050 150.820 125.380 152.430 ;
        RECT 122.810 150.400 123.510 150.570 ;
        RECT 124.180 150.400 124.880 150.570 ;
        RECT 122.310 148.540 122.640 150.150 ;
        RECT 123.680 148.540 124.010 150.150 ;
        RECT 125.050 148.540 125.380 150.150 ;
        RECT 122.810 148.120 123.510 148.290 ;
        RECT 124.180 148.120 124.880 148.290 ;
        RECT 122.310 146.260 122.640 147.870 ;
        RECT 123.680 146.260 124.010 147.870 ;
        RECT 125.050 146.260 125.380 147.870 ;
        RECT 122.810 145.840 123.510 146.010 ;
        RECT 124.180 145.840 124.880 146.010 ;
        RECT 122.310 143.980 122.640 145.590 ;
        RECT 123.680 143.980 124.010 145.590 ;
        RECT 125.050 143.980 125.380 145.590 ;
        RECT 122.810 143.560 123.510 143.730 ;
        RECT 124.180 143.560 124.880 143.730 ;
        RECT 122.310 141.700 122.640 143.310 ;
        RECT 123.680 141.700 124.010 143.310 ;
        RECT 125.050 141.700 125.380 143.310 ;
        RECT 122.810 141.280 123.510 141.450 ;
        RECT 124.180 141.280 124.880 141.450 ;
        RECT 122.310 139.420 122.640 141.030 ;
        RECT 123.680 139.420 124.010 141.030 ;
        RECT 125.050 139.420 125.380 141.030 ;
        RECT 122.810 139.000 123.510 139.170 ;
        RECT 124.180 139.000 124.880 139.170 ;
        RECT 122.310 137.140 122.640 138.750 ;
        RECT 123.680 137.140 124.010 138.750 ;
        RECT 125.050 137.140 125.380 138.750 ;
        RECT 122.810 136.720 123.510 136.890 ;
        RECT 124.180 136.720 124.880 136.890 ;
        RECT 122.310 134.860 122.640 136.470 ;
        RECT 123.680 134.860 124.010 136.470 ;
        RECT 125.050 134.860 125.380 136.470 ;
        RECT 122.810 134.440 123.510 134.610 ;
        RECT 124.180 134.440 124.880 134.610 ;
        RECT 122.310 132.580 122.640 134.190 ;
        RECT 123.680 132.580 124.010 134.190 ;
        RECT 125.050 132.580 125.380 134.190 ;
        RECT 122.810 132.160 123.510 132.330 ;
        RECT 124.180 132.160 124.880 132.330 ;
        RECT 122.310 130.300 122.640 131.910 ;
        RECT 123.680 130.300 124.010 131.910 ;
        RECT 125.050 130.300 125.380 131.910 ;
        RECT 122.810 129.880 123.510 130.050 ;
        RECT 124.180 129.880 124.880 130.050 ;
        RECT 122.310 128.020 122.640 129.630 ;
        RECT 123.680 128.020 124.010 129.630 ;
        RECT 125.050 128.020 125.380 129.630 ;
        RECT 122.810 127.600 123.510 127.770 ;
        RECT 124.180 127.600 124.880 127.770 ;
        RECT 122.310 125.740 122.640 127.350 ;
        RECT 123.680 125.740 124.010 127.350 ;
        RECT 125.050 125.740 125.380 127.350 ;
        RECT 122.810 125.320 123.510 125.490 ;
        RECT 124.180 125.320 124.880 125.490 ;
        RECT 122.310 123.460 122.640 125.070 ;
        RECT 123.680 123.460 124.010 125.070 ;
        RECT 125.050 123.460 125.380 125.070 ;
        RECT 122.810 123.040 123.510 123.210 ;
        RECT 124.180 123.040 124.880 123.210 ;
        RECT 122.310 121.180 122.640 122.790 ;
        RECT 123.680 121.180 124.010 122.790 ;
        RECT 125.050 121.180 125.380 122.790 ;
        RECT 122.810 120.760 123.510 120.930 ;
        RECT 124.180 120.760 124.880 120.930 ;
        RECT 122.310 118.900 122.640 120.510 ;
        RECT 123.680 118.900 124.010 120.510 ;
        RECT 125.050 118.900 125.380 120.510 ;
        RECT 122.810 118.480 123.510 118.650 ;
        RECT 124.180 118.480 124.880 118.650 ;
        RECT 122.310 116.620 122.640 118.230 ;
        RECT 123.680 116.620 124.010 118.230 ;
        RECT 125.050 116.620 125.380 118.230 ;
        RECT 122.810 116.200 123.510 116.370 ;
        RECT 124.180 116.200 124.880 116.370 ;
        RECT 122.310 114.340 122.640 115.950 ;
        RECT 123.680 114.340 124.010 115.950 ;
        RECT 125.050 114.340 125.380 115.950 ;
        RECT 122.810 113.920 123.510 114.090 ;
        RECT 124.180 113.920 124.880 114.090 ;
        RECT 122.310 112.060 122.640 113.670 ;
        RECT 123.680 112.060 124.010 113.670 ;
        RECT 125.050 112.060 125.380 113.670 ;
        RECT 122.810 111.640 123.510 111.810 ;
        RECT 124.180 111.640 124.880 111.810 ;
        RECT 122.310 109.780 122.640 111.390 ;
        RECT 123.680 109.780 124.010 111.390 ;
        RECT 125.050 109.780 125.380 111.390 ;
        RECT 122.810 109.360 123.510 109.530 ;
        RECT 124.180 109.360 124.880 109.530 ;
        RECT 122.310 107.500 122.640 109.110 ;
        RECT 123.680 107.500 124.010 109.110 ;
        RECT 125.050 107.500 125.380 109.110 ;
        RECT 122.810 107.080 123.510 107.250 ;
        RECT 124.180 107.080 124.880 107.250 ;
        RECT 122.310 105.220 122.640 106.830 ;
        RECT 123.680 105.220 124.010 106.830 ;
        RECT 125.050 105.220 125.380 106.830 ;
        RECT 122.810 104.800 123.510 104.970 ;
        RECT 124.180 104.800 124.880 104.970 ;
        RECT 122.310 102.940 122.640 104.550 ;
        RECT 123.680 102.940 124.010 104.550 ;
        RECT 125.050 102.940 125.380 104.550 ;
        RECT 122.810 102.520 123.510 102.690 ;
        RECT 124.180 102.520 124.880 102.690 ;
        RECT 122.310 100.660 122.640 102.270 ;
        RECT 123.680 100.660 124.010 102.270 ;
        RECT 125.050 100.660 125.380 102.270 ;
        RECT 122.810 100.240 123.510 100.410 ;
        RECT 124.180 100.240 124.880 100.410 ;
        RECT 122.310 98.380 122.640 99.990 ;
        RECT 123.680 98.380 124.010 99.990 ;
        RECT 125.050 98.380 125.380 99.990 ;
        RECT 122.810 97.960 123.510 98.130 ;
        RECT 124.180 97.960 124.880 98.130 ;
        RECT 122.310 96.100 122.640 97.710 ;
        RECT 123.680 96.100 124.010 97.710 ;
        RECT 125.050 96.100 125.380 97.710 ;
        RECT 122.810 95.680 123.510 95.850 ;
        RECT 124.180 95.680 124.880 95.850 ;
        RECT 122.310 93.820 122.640 95.430 ;
        RECT 123.680 93.820 124.010 95.430 ;
        RECT 125.050 93.820 125.380 95.430 ;
        RECT 122.810 93.400 123.510 93.570 ;
        RECT 124.180 93.400 124.880 93.570 ;
        RECT 122.310 91.540 122.640 93.150 ;
        RECT 123.680 91.540 124.010 93.150 ;
        RECT 125.050 91.540 125.380 93.150 ;
        RECT 122.810 91.120 123.510 91.290 ;
        RECT 124.180 91.120 124.880 91.290 ;
        RECT 122.310 89.260 122.640 90.870 ;
        RECT 125.050 89.260 125.380 90.870 ;
        RECT 122.810 88.840 123.510 89.010 ;
        RECT 124.180 88.840 124.880 89.010 ;
        RECT 122.310 86.980 122.640 88.590 ;
        RECT 125.050 86.980 125.380 88.590 ;
        RECT 122.810 86.560 123.510 86.730 ;
        RECT 124.180 86.560 124.880 86.730 ;
        RECT 122.310 84.700 122.640 86.310 ;
        RECT 125.050 84.700 125.380 86.310 ;
        RECT 122.810 84.280 123.510 84.450 ;
        RECT 124.180 84.280 124.880 84.450 ;
        RECT 122.310 82.420 122.640 84.030 ;
        RECT 125.050 82.420 125.380 84.030 ;
        RECT 122.810 82.000 123.510 82.170 ;
        RECT 124.180 82.000 124.880 82.170 ;
        RECT 122.310 80.140 122.640 81.750 ;
        RECT 125.050 80.140 125.380 81.750 ;
        RECT 122.810 79.720 123.510 79.890 ;
        RECT 124.180 79.720 124.880 79.890 ;
        RECT 122.310 77.860 122.640 79.470 ;
        RECT 123.680 77.860 124.010 79.470 ;
        RECT 125.050 77.860 125.380 79.470 ;
        RECT 122.810 77.440 123.510 77.610 ;
        RECT 124.180 77.440 124.880 77.610 ;
        RECT 125.680 76.980 125.850 164.710 ;
        RECT 121.840 76.810 125.850 76.980 ;
        RECT 118.195 75.580 121.135 75.750 ;
        RECT 114.925 75.405 117.565 75.575 ;
        RECT 108.635 63.090 114.015 63.260 ;
        RECT 114.775 70.630 117.415 70.800 ;
        RECT 114.775 60.340 114.945 70.630 ;
        RECT 115.745 69.960 116.445 70.130 ;
        RECT 116.615 68.100 116.945 69.710 ;
        RECT 115.745 67.680 116.445 67.850 ;
        RECT 115.245 65.820 115.575 67.430 ;
        RECT 115.745 65.400 116.445 65.570 ;
        RECT 115.245 63.540 115.575 65.150 ;
        RECT 115.745 63.120 116.445 63.290 ;
        RECT 116.615 61.260 116.945 62.870 ;
        RECT 115.745 60.840 116.445 61.010 ;
        RECT 117.245 60.340 117.415 70.630 ;
        RECT 118.470 70.350 123.825 70.520 ;
        RECT 118.470 65.740 118.640 70.350 ;
        RECT 119.440 69.680 120.140 69.850 ;
        RECT 122.155 69.680 122.855 69.850 ;
        RECT 118.940 69.250 119.270 69.420 ;
        RECT 119.440 69.250 120.140 69.420 ;
        RECT 121.655 69.250 121.985 69.420 ;
        RECT 122.155 69.250 122.855 69.420 ;
        RECT 119.440 68.820 120.140 68.990 ;
        RECT 122.155 68.820 122.855 68.990 ;
        RECT 119.440 68.390 120.140 68.560 ;
        RECT 120.310 68.390 120.640 68.560 ;
        RECT 122.155 68.390 122.855 68.560 ;
        RECT 123.025 68.390 123.355 68.560 ;
        RECT 119.440 67.960 120.140 68.130 ;
        RECT 122.155 67.960 122.855 68.130 ;
        RECT 119.440 67.530 120.140 67.700 ;
        RECT 120.310 67.530 120.640 67.700 ;
        RECT 122.155 67.530 122.855 67.700 ;
        RECT 123.025 67.530 123.355 67.700 ;
        RECT 119.440 67.100 120.140 67.270 ;
        RECT 122.155 67.100 122.855 67.270 ;
        RECT 118.940 66.670 119.270 66.840 ;
        RECT 119.440 66.670 120.140 66.840 ;
        RECT 121.655 66.670 121.985 66.840 ;
        RECT 122.155 66.670 122.855 66.840 ;
        RECT 119.440 66.240 120.140 66.410 ;
        RECT 122.155 66.240 122.855 66.410 ;
        RECT 123.655 65.740 123.825 70.350 ;
        RECT 118.470 65.570 123.825 65.740 ;
        RECT 124.455 70.310 127.095 70.480 ;
        RECT 118.470 65.060 123.825 65.230 ;
        RECT 118.470 60.530 118.640 65.060 ;
        RECT 119.440 64.430 120.140 64.600 ;
        RECT 122.155 64.430 122.855 64.600 ;
        RECT 118.940 64.000 119.270 64.170 ;
        RECT 119.440 64.000 120.140 64.170 ;
        RECT 121.655 64.000 121.985 64.170 ;
        RECT 122.155 64.000 122.855 64.170 ;
        RECT 119.440 63.570 120.140 63.740 ;
        RECT 122.155 63.570 122.855 63.740 ;
        RECT 119.440 63.140 120.140 63.310 ;
        RECT 120.310 63.140 120.640 63.310 ;
        RECT 122.155 63.140 122.855 63.310 ;
        RECT 123.025 63.140 123.355 63.310 ;
        RECT 119.440 62.710 120.140 62.880 ;
        RECT 122.155 62.710 122.855 62.880 ;
        RECT 119.440 62.280 120.140 62.450 ;
        RECT 120.310 62.280 120.640 62.450 ;
        RECT 122.155 62.280 122.855 62.450 ;
        RECT 123.025 62.280 123.355 62.450 ;
        RECT 119.440 61.850 120.140 62.020 ;
        RECT 122.155 61.850 122.855 62.020 ;
        RECT 118.940 61.420 119.270 61.590 ;
        RECT 119.440 61.420 120.140 61.590 ;
        RECT 121.655 61.420 121.985 61.590 ;
        RECT 122.155 61.420 122.855 61.590 ;
        RECT 119.440 60.990 120.140 61.160 ;
        RECT 122.155 60.990 122.855 61.160 ;
        RECT 123.655 60.530 123.825 65.060 ;
        RECT 118.470 60.360 123.825 60.530 ;
        RECT 124.455 60.620 124.625 70.310 ;
        RECT 125.425 69.680 126.125 69.850 ;
        RECT 124.925 69.250 125.255 69.420 ;
        RECT 125.425 69.250 126.125 69.420 ;
        RECT 125.425 68.820 126.125 68.990 ;
        RECT 124.925 68.390 125.255 68.560 ;
        RECT 125.425 68.390 126.125 68.560 ;
        RECT 125.425 67.960 126.125 68.130 ;
        RECT 124.925 67.530 125.255 67.700 ;
        RECT 125.425 67.530 126.125 67.700 ;
        RECT 125.425 67.100 126.125 67.270 ;
        RECT 124.925 66.670 125.255 66.840 ;
        RECT 125.425 66.670 126.125 66.840 ;
        RECT 125.425 66.240 126.125 66.410 ;
        RECT 125.425 65.810 126.125 65.980 ;
        RECT 126.295 65.810 126.625 65.980 ;
        RECT 125.425 65.380 126.125 65.550 ;
        RECT 125.425 64.950 126.125 65.120 ;
        RECT 126.295 64.950 126.625 65.120 ;
        RECT 125.425 64.520 126.125 64.690 ;
        RECT 124.925 64.090 125.255 64.260 ;
        RECT 125.425 64.090 126.125 64.260 ;
        RECT 125.425 63.660 126.125 63.830 ;
        RECT 124.925 63.230 125.255 63.400 ;
        RECT 125.425 63.230 126.125 63.400 ;
        RECT 125.425 62.800 126.125 62.970 ;
        RECT 124.925 62.370 125.255 62.540 ;
        RECT 125.425 62.370 126.125 62.540 ;
        RECT 125.425 61.940 126.125 62.110 ;
        RECT 124.925 61.510 125.255 61.680 ;
        RECT 125.425 61.510 126.125 61.680 ;
        RECT 125.425 61.080 126.125 61.250 ;
        RECT 126.925 60.620 127.095 70.310 ;
        RECT 124.455 60.450 127.095 60.620 ;
        RECT 114.775 60.170 117.415 60.340 ;
      LAYER mcon ;
        RECT 107.890 173.900 108.060 174.070 ;
        RECT 108.250 173.900 108.420 174.070 ;
        RECT 108.610 173.900 108.780 174.070 ;
        RECT 108.970 173.900 109.140 174.070 ;
        RECT 109.330 173.900 109.500 174.070 ;
        RECT 109.690 173.900 109.860 174.070 ;
        RECT 111.185 173.900 111.355 174.070 ;
        RECT 111.545 173.900 111.715 174.070 ;
        RECT 111.905 173.900 112.075 174.070 ;
        RECT 112.265 173.900 112.435 174.070 ;
        RECT 112.625 173.900 112.795 174.070 ;
        RECT 112.985 173.900 113.155 174.070 ;
        RECT 113.345 173.900 113.515 174.070 ;
        RECT 113.705 173.900 113.875 174.070 ;
        RECT 107.590 173.550 107.760 173.720 ;
        RECT 114.005 173.550 114.175 173.720 ;
        RECT 107.590 173.190 107.760 173.360 ;
        RECT 108.430 173.230 108.600 173.400 ;
        RECT 108.790 173.230 108.960 173.400 ;
        RECT 111.740 173.230 111.910 173.400 ;
        RECT 112.100 173.230 112.270 173.400 ;
        RECT 112.460 173.230 112.630 173.400 ;
        RECT 112.820 173.230 112.990 173.400 ;
        RECT 113.180 173.230 113.350 173.400 ;
        RECT 114.005 173.190 114.175 173.360 ;
        RECT 107.590 172.830 107.760 173.000 ;
        RECT 109.445 172.980 109.615 173.150 ;
        RECT 108.430 172.800 108.600 172.970 ;
        RECT 108.790 172.800 108.960 172.970 ;
        RECT 107.590 172.470 107.760 172.640 ;
        RECT 109.445 172.620 109.615 172.790 ;
        RECT 111.125 172.980 111.295 173.150 ;
        RECT 111.740 172.800 111.910 172.970 ;
        RECT 112.100 172.800 112.270 172.970 ;
        RECT 112.460 172.800 112.630 172.970 ;
        RECT 112.820 172.800 112.990 172.970 ;
        RECT 113.180 172.800 113.350 172.970 ;
        RECT 114.005 172.830 114.175 173.000 ;
        RECT 111.125 172.620 111.295 172.790 ;
        RECT 108.430 172.370 108.600 172.540 ;
        RECT 108.790 172.370 108.960 172.540 ;
        RECT 111.740 172.370 111.910 172.540 ;
        RECT 112.100 172.370 112.270 172.540 ;
        RECT 112.460 172.370 112.630 172.540 ;
        RECT 112.820 172.370 112.990 172.540 ;
        RECT 113.180 172.370 113.350 172.540 ;
        RECT 114.005 172.470 114.175 172.640 ;
        RECT 107.590 172.110 107.760 172.280 ;
        RECT 109.445 172.120 109.615 172.290 ;
        RECT 108.430 171.940 108.600 172.110 ;
        RECT 108.790 171.940 108.960 172.110 ;
        RECT 107.590 171.750 107.760 171.920 ;
        RECT 109.445 171.760 109.615 171.930 ;
        RECT 111.125 172.120 111.295 172.290 ;
        RECT 114.005 172.110 114.175 172.280 ;
        RECT 111.740 171.940 111.910 172.110 ;
        RECT 112.100 171.940 112.270 172.110 ;
        RECT 112.460 171.940 112.630 172.110 ;
        RECT 112.820 171.940 112.990 172.110 ;
        RECT 113.180 171.940 113.350 172.110 ;
        RECT 111.125 171.760 111.295 171.930 ;
        RECT 114.005 171.750 114.175 171.920 ;
        RECT 107.590 171.390 107.760 171.560 ;
        RECT 108.430 171.510 108.600 171.680 ;
        RECT 108.790 171.510 108.960 171.680 ;
        RECT 111.740 171.510 111.910 171.680 ;
        RECT 112.100 171.510 112.270 171.680 ;
        RECT 112.460 171.510 112.630 171.680 ;
        RECT 112.820 171.510 112.990 171.680 ;
        RECT 113.180 171.510 113.350 171.680 ;
        RECT 109.445 171.260 109.615 171.430 ;
        RECT 107.590 171.030 107.760 171.200 ;
        RECT 108.430 171.080 108.600 171.250 ;
        RECT 108.790 171.080 108.960 171.250 ;
        RECT 109.445 170.900 109.615 171.070 ;
        RECT 111.125 171.260 111.295 171.430 ;
        RECT 114.005 171.390 114.175 171.560 ;
        RECT 111.740 171.080 111.910 171.250 ;
        RECT 112.100 171.080 112.270 171.250 ;
        RECT 112.460 171.080 112.630 171.250 ;
        RECT 112.820 171.080 112.990 171.250 ;
        RECT 113.180 171.080 113.350 171.250 ;
        RECT 111.125 170.900 111.295 171.070 ;
        RECT 114.005 171.030 114.175 171.200 ;
        RECT 107.590 170.670 107.760 170.840 ;
        RECT 108.430 170.650 108.600 170.820 ;
        RECT 108.790 170.650 108.960 170.820 ;
        RECT 111.740 170.650 111.910 170.820 ;
        RECT 112.100 170.650 112.270 170.820 ;
        RECT 112.460 170.650 112.630 170.820 ;
        RECT 112.820 170.650 112.990 170.820 ;
        RECT 113.180 170.650 113.350 170.820 ;
        RECT 114.005 170.670 114.175 170.840 ;
        RECT 107.590 170.310 107.760 170.480 ;
        RECT 109.445 170.400 109.615 170.570 ;
        RECT 108.430 170.220 108.600 170.390 ;
        RECT 108.790 170.220 108.960 170.390 ;
        RECT 107.590 169.950 107.760 170.120 ;
        RECT 109.445 170.040 109.615 170.210 ;
        RECT 111.125 170.400 111.295 170.570 ;
        RECT 111.740 170.220 111.910 170.390 ;
        RECT 112.100 170.220 112.270 170.390 ;
        RECT 112.460 170.220 112.630 170.390 ;
        RECT 112.820 170.220 112.990 170.390 ;
        RECT 113.180 170.220 113.350 170.390 ;
        RECT 114.005 170.310 114.175 170.480 ;
        RECT 111.125 170.040 111.295 170.210 ;
        RECT 108.430 169.790 108.600 169.960 ;
        RECT 108.790 169.790 108.960 169.960 ;
        RECT 111.740 169.790 111.910 169.960 ;
        RECT 112.100 169.790 112.270 169.960 ;
        RECT 112.460 169.790 112.630 169.960 ;
        RECT 112.820 169.790 112.990 169.960 ;
        RECT 113.180 169.790 113.350 169.960 ;
        RECT 114.005 169.950 114.175 170.120 ;
        RECT 107.590 169.590 107.760 169.760 ;
        RECT 114.005 169.590 114.175 169.760 ;
        RECT 107.890 169.120 108.060 169.290 ;
        RECT 108.250 169.120 108.420 169.290 ;
        RECT 108.610 169.120 108.780 169.290 ;
        RECT 108.970 169.120 109.140 169.290 ;
        RECT 109.330 169.120 109.500 169.290 ;
        RECT 109.690 169.120 109.860 169.290 ;
        RECT 111.185 169.120 111.355 169.290 ;
        RECT 111.545 169.120 111.715 169.290 ;
        RECT 111.905 169.120 112.075 169.290 ;
        RECT 112.265 169.120 112.435 169.290 ;
        RECT 112.625 169.120 112.795 169.290 ;
        RECT 112.985 169.120 113.155 169.290 ;
        RECT 113.345 169.120 113.515 169.290 ;
        RECT 113.705 169.120 113.875 169.290 ;
        RECT 108.635 164.690 108.805 164.860 ;
        RECT 109.105 164.750 109.275 164.920 ;
        RECT 109.465 164.750 109.635 164.920 ;
        RECT 109.825 164.750 109.995 164.920 ;
        RECT 110.185 164.750 110.355 164.920 ;
        RECT 110.545 164.750 110.715 164.920 ;
        RECT 110.905 164.750 111.075 164.920 ;
        RECT 111.265 164.750 111.435 164.920 ;
        RECT 111.625 164.750 111.795 164.920 ;
        RECT 111.985 164.750 112.155 164.920 ;
        RECT 112.345 164.750 112.515 164.920 ;
        RECT 112.705 164.750 112.875 164.920 ;
        RECT 113.065 164.750 113.235 164.920 ;
        RECT 113.425 164.750 113.595 164.920 ;
        RECT 113.785 164.750 113.955 164.920 ;
        RECT 108.635 164.330 108.805 164.500 ;
        RECT 113.845 164.310 114.015 164.480 ;
        RECT 108.635 163.970 108.805 164.140 ;
        RECT 109.690 164.080 109.860 164.250 ;
        RECT 110.050 164.080 110.220 164.250 ;
        RECT 111.060 164.080 111.230 164.250 ;
        RECT 111.420 164.080 111.590 164.250 ;
        RECT 112.430 164.080 112.600 164.250 ;
        RECT 112.790 164.080 112.960 164.250 ;
        RECT 113.845 163.950 114.015 164.120 ;
        RECT 108.635 163.610 108.805 163.780 ;
        RECT 108.635 163.250 108.805 163.420 ;
        RECT 108.635 162.890 108.805 163.060 ;
        RECT 108.635 162.530 108.805 162.700 ;
        RECT 108.635 162.170 108.805 162.340 ;
        RECT 110.555 163.660 110.725 163.830 ;
        RECT 110.555 163.300 110.725 163.470 ;
        RECT 110.555 162.940 110.725 163.110 ;
        RECT 110.555 162.580 110.725 162.750 ;
        RECT 110.555 162.220 110.725 162.390 ;
        RECT 111.925 163.660 112.095 163.830 ;
        RECT 111.925 163.300 112.095 163.470 ;
        RECT 111.925 162.940 112.095 163.110 ;
        RECT 111.925 162.580 112.095 162.750 ;
        RECT 111.925 162.220 112.095 162.390 ;
        RECT 113.845 163.590 114.015 163.760 ;
        RECT 113.845 163.230 114.015 163.400 ;
        RECT 113.845 162.870 114.015 163.040 ;
        RECT 113.845 162.510 114.015 162.680 ;
        RECT 108.635 161.810 108.805 161.980 ;
        RECT 113.845 162.150 114.015 162.320 ;
        RECT 109.690 161.800 109.860 161.970 ;
        RECT 110.050 161.800 110.220 161.970 ;
        RECT 111.060 161.800 111.230 161.970 ;
        RECT 111.420 161.800 111.590 161.970 ;
        RECT 112.430 161.800 112.600 161.970 ;
        RECT 112.790 161.800 112.960 161.970 ;
        RECT 108.635 161.450 108.805 161.620 ;
        RECT 113.845 161.790 114.015 161.960 ;
        RECT 108.635 161.090 108.805 161.260 ;
        RECT 108.635 160.730 108.805 160.900 ;
        RECT 108.635 160.370 108.805 160.540 ;
        RECT 108.635 160.010 108.805 160.180 ;
        RECT 110.555 161.380 110.725 161.550 ;
        RECT 110.555 161.020 110.725 161.190 ;
        RECT 110.555 160.660 110.725 160.830 ;
        RECT 110.555 160.300 110.725 160.470 ;
        RECT 110.555 159.940 110.725 160.110 ;
        RECT 111.925 161.380 112.095 161.550 ;
        RECT 111.925 161.020 112.095 161.190 ;
        RECT 111.925 160.660 112.095 160.830 ;
        RECT 111.925 160.300 112.095 160.470 ;
        RECT 111.925 159.940 112.095 160.110 ;
        RECT 113.845 161.430 114.015 161.600 ;
        RECT 113.845 161.070 114.015 161.240 ;
        RECT 113.845 160.710 114.015 160.880 ;
        RECT 113.845 160.350 114.015 160.520 ;
        RECT 113.845 159.990 114.015 160.160 ;
        RECT 108.635 159.650 108.805 159.820 ;
        RECT 109.690 159.520 109.860 159.690 ;
        RECT 110.050 159.520 110.220 159.690 ;
        RECT 111.060 159.520 111.230 159.690 ;
        RECT 111.420 159.520 111.590 159.690 ;
        RECT 112.430 159.520 112.600 159.690 ;
        RECT 112.790 159.520 112.960 159.690 ;
        RECT 113.845 159.630 114.015 159.800 ;
        RECT 108.635 159.290 108.805 159.460 ;
        RECT 113.845 159.270 114.015 159.440 ;
        RECT 108.635 158.930 108.805 159.100 ;
        RECT 108.635 158.570 108.805 158.740 ;
        RECT 108.635 158.210 108.805 158.380 ;
        RECT 108.635 157.850 108.805 158.020 ;
        RECT 110.555 159.100 110.725 159.270 ;
        RECT 110.555 158.740 110.725 158.910 ;
        RECT 110.555 158.380 110.725 158.550 ;
        RECT 110.555 158.020 110.725 158.190 ;
        RECT 110.555 157.660 110.725 157.830 ;
        RECT 111.925 159.100 112.095 159.270 ;
        RECT 111.925 158.740 112.095 158.910 ;
        RECT 111.925 158.380 112.095 158.550 ;
        RECT 111.925 158.020 112.095 158.190 ;
        RECT 111.925 157.660 112.095 157.830 ;
        RECT 113.845 158.910 114.015 159.080 ;
        RECT 113.845 158.550 114.015 158.720 ;
        RECT 113.845 158.190 114.015 158.360 ;
        RECT 113.845 157.830 114.015 158.000 ;
        RECT 108.635 157.490 108.805 157.660 ;
        RECT 113.845 157.470 114.015 157.640 ;
        RECT 108.635 157.130 108.805 157.300 ;
        RECT 109.690 157.240 109.860 157.410 ;
        RECT 110.050 157.240 110.220 157.410 ;
        RECT 111.060 157.240 111.230 157.410 ;
        RECT 111.420 157.240 111.590 157.410 ;
        RECT 112.430 157.240 112.600 157.410 ;
        RECT 112.790 157.240 112.960 157.410 ;
        RECT 113.845 157.110 114.015 157.280 ;
        RECT 108.635 156.770 108.805 156.940 ;
        RECT 108.635 156.410 108.805 156.580 ;
        RECT 108.635 156.050 108.805 156.220 ;
        RECT 108.635 155.690 108.805 155.860 ;
        RECT 108.635 155.330 108.805 155.500 ;
        RECT 110.555 156.820 110.725 156.990 ;
        RECT 110.555 156.460 110.725 156.630 ;
        RECT 110.555 156.100 110.725 156.270 ;
        RECT 110.555 155.740 110.725 155.910 ;
        RECT 110.555 155.380 110.725 155.550 ;
        RECT 111.925 156.820 112.095 156.990 ;
        RECT 111.925 156.460 112.095 156.630 ;
        RECT 111.925 156.100 112.095 156.270 ;
        RECT 111.925 155.740 112.095 155.910 ;
        RECT 111.925 155.380 112.095 155.550 ;
        RECT 113.845 156.750 114.015 156.920 ;
        RECT 113.845 156.390 114.015 156.560 ;
        RECT 113.845 156.030 114.015 156.200 ;
        RECT 113.845 155.670 114.015 155.840 ;
        RECT 108.635 154.970 108.805 155.140 ;
        RECT 113.845 155.310 114.015 155.480 ;
        RECT 109.690 154.960 109.860 155.130 ;
        RECT 110.050 154.960 110.220 155.130 ;
        RECT 111.060 154.960 111.230 155.130 ;
        RECT 111.420 154.960 111.590 155.130 ;
        RECT 112.430 154.960 112.600 155.130 ;
        RECT 112.790 154.960 112.960 155.130 ;
        RECT 108.635 154.610 108.805 154.780 ;
        RECT 113.845 154.950 114.015 155.120 ;
        RECT 108.635 154.250 108.805 154.420 ;
        RECT 108.635 153.890 108.805 154.060 ;
        RECT 108.635 153.530 108.805 153.700 ;
        RECT 108.635 153.170 108.805 153.340 ;
        RECT 110.555 154.540 110.725 154.710 ;
        RECT 110.555 154.180 110.725 154.350 ;
        RECT 110.555 153.820 110.725 153.990 ;
        RECT 110.555 153.460 110.725 153.630 ;
        RECT 110.555 153.100 110.725 153.270 ;
        RECT 111.925 154.540 112.095 154.710 ;
        RECT 111.925 154.180 112.095 154.350 ;
        RECT 111.925 153.820 112.095 153.990 ;
        RECT 111.925 153.460 112.095 153.630 ;
        RECT 111.925 153.100 112.095 153.270 ;
        RECT 113.845 154.590 114.015 154.760 ;
        RECT 113.845 154.230 114.015 154.400 ;
        RECT 113.845 153.870 114.015 154.040 ;
        RECT 113.845 153.510 114.015 153.680 ;
        RECT 113.845 153.150 114.015 153.320 ;
        RECT 108.635 152.810 108.805 152.980 ;
        RECT 109.690 152.680 109.860 152.850 ;
        RECT 110.050 152.680 110.220 152.850 ;
        RECT 111.060 152.680 111.230 152.850 ;
        RECT 111.420 152.680 111.590 152.850 ;
        RECT 112.430 152.680 112.600 152.850 ;
        RECT 112.790 152.680 112.960 152.850 ;
        RECT 113.845 152.790 114.015 152.960 ;
        RECT 108.635 152.450 108.805 152.620 ;
        RECT 113.845 152.430 114.015 152.600 ;
        RECT 108.635 152.090 108.805 152.260 ;
        RECT 108.635 151.730 108.805 151.900 ;
        RECT 56.480 151.500 56.650 151.670 ;
        RECT 56.840 151.500 57.010 151.670 ;
        RECT 57.200 151.500 57.370 151.670 ;
        RECT 57.560 151.500 57.730 151.670 ;
        RECT 57.920 151.500 58.090 151.670 ;
        RECT 58.280 151.500 58.450 151.670 ;
        RECT 58.640 151.500 58.810 151.670 ;
        RECT 59.000 151.500 59.170 151.670 ;
        RECT 59.360 151.500 59.530 151.670 ;
        RECT 59.720 151.500 59.890 151.670 ;
        RECT 60.080 151.500 60.250 151.670 ;
        RECT 60.440 151.500 60.610 151.670 ;
        RECT 60.800 151.500 60.970 151.670 ;
        RECT 61.160 151.500 61.330 151.670 ;
        RECT 61.520 151.500 61.690 151.670 ;
        RECT 61.880 151.500 62.050 151.670 ;
        RECT 62.240 151.500 62.410 151.670 ;
        RECT 56.180 151.150 56.350 151.320 ;
        RECT 62.540 151.150 62.710 151.320 ;
        RECT 56.180 150.790 56.350 150.960 ;
        RECT 60.975 150.830 61.145 151.000 ;
        RECT 61.335 150.830 61.505 151.000 ;
        RECT 56.180 150.430 56.350 150.600 ;
        RECT 62.540 150.790 62.710 150.960 ;
        RECT 56.180 150.070 56.350 150.240 ;
        RECT 56.180 149.710 56.350 149.880 ;
        RECT 60.320 150.410 60.490 150.580 ;
        RECT 62.540 150.430 62.710 150.600 ;
        RECT 60.320 150.050 60.490 150.220 ;
        RECT 60.975 150.050 61.145 150.220 ;
        RECT 61.335 150.050 61.505 150.220 ;
        RECT 62.540 150.070 62.710 150.240 ;
        RECT 60.320 149.690 60.490 149.860 ;
        RECT 62.540 149.710 62.710 149.880 ;
        RECT 56.180 149.350 56.350 149.520 ;
        RECT 60.975 149.270 61.145 149.440 ;
        RECT 61.335 149.270 61.505 149.440 ;
        RECT 62.540 149.350 62.710 149.520 ;
        RECT 56.180 148.990 56.350 149.160 ;
        RECT 56.180 148.630 56.350 148.800 ;
        RECT 56.180 148.270 56.350 148.440 ;
        RECT 56.180 147.910 56.350 148.080 ;
        RECT 56.180 147.550 56.350 147.720 ;
        RECT 61.990 148.850 62.160 149.020 ;
        RECT 61.990 148.490 62.160 148.660 ;
        RECT 61.990 148.130 62.160 148.300 ;
        RECT 61.990 147.770 62.160 147.940 ;
        RECT 61.990 147.410 62.160 147.580 ;
        RECT 62.540 148.990 62.710 149.160 ;
        RECT 62.540 148.630 62.710 148.800 ;
        RECT 62.540 148.270 62.710 148.440 ;
        RECT 62.540 147.910 62.710 148.080 ;
        RECT 62.540 147.550 62.710 147.720 ;
        RECT 56.180 147.190 56.350 147.360 ;
        RECT 62.540 147.190 62.710 147.360 ;
        RECT 56.180 146.830 56.350 147.000 ;
        RECT 60.975 146.990 61.145 147.160 ;
        RECT 61.335 146.990 61.505 147.160 ;
        RECT 62.540 146.830 62.710 147.000 ;
        RECT 56.180 146.470 56.350 146.640 ;
        RECT 56.180 146.110 56.350 146.280 ;
        RECT 56.180 145.750 56.350 145.920 ;
        RECT 56.180 145.390 56.350 145.560 ;
        RECT 56.180 145.030 56.350 145.200 ;
        RECT 61.990 146.570 62.160 146.740 ;
        RECT 61.990 146.210 62.160 146.380 ;
        RECT 61.990 145.850 62.160 146.020 ;
        RECT 61.990 145.490 62.160 145.660 ;
        RECT 61.990 145.130 62.160 145.300 ;
        RECT 62.540 146.470 62.710 146.640 ;
        RECT 62.540 146.110 62.710 146.280 ;
        RECT 62.540 145.750 62.710 145.920 ;
        RECT 62.540 145.390 62.710 145.560 ;
        RECT 62.540 145.030 62.710 145.200 ;
        RECT 56.180 144.670 56.350 144.840 ;
        RECT 60.975 144.710 61.145 144.880 ;
        RECT 61.335 144.710 61.505 144.880 ;
        RECT 56.180 144.310 56.350 144.480 ;
        RECT 62.540 144.670 62.710 144.840 ;
        RECT 56.180 143.950 56.350 144.120 ;
        RECT 56.180 143.590 56.350 143.760 ;
        RECT 60.320 144.290 60.490 144.460 ;
        RECT 62.540 144.310 62.710 144.480 ;
        RECT 60.320 143.930 60.490 144.100 ;
        RECT 60.975 143.930 61.145 144.100 ;
        RECT 61.335 143.930 61.505 144.100 ;
        RECT 62.540 143.950 62.710 144.120 ;
        RECT 60.320 143.570 60.490 143.740 ;
        RECT 62.540 143.590 62.710 143.760 ;
        RECT 56.180 143.230 56.350 143.400 ;
        RECT 60.975 143.150 61.145 143.320 ;
        RECT 61.335 143.150 61.505 143.320 ;
        RECT 62.540 143.230 62.710 143.400 ;
        RECT 56.180 142.870 56.350 143.040 ;
        RECT 56.180 142.510 56.350 142.680 ;
        RECT 56.180 142.150 56.350 142.320 ;
        RECT 60.320 142.730 60.490 142.900 ;
        RECT 62.540 142.870 62.710 143.040 ;
        RECT 60.320 142.370 60.490 142.540 ;
        RECT 60.975 142.370 61.145 142.540 ;
        RECT 61.335 142.370 61.505 142.540 ;
        RECT 62.540 142.510 62.710 142.680 ;
        RECT 60.320 142.010 60.490 142.180 ;
        RECT 64.965 151.500 65.135 151.670 ;
        RECT 65.325 151.500 65.495 151.670 ;
        RECT 65.685 151.500 65.855 151.670 ;
        RECT 66.045 151.500 66.215 151.670 ;
        RECT 66.405 151.500 66.575 151.670 ;
        RECT 64.435 151.150 64.605 151.320 ;
        RECT 66.705 151.150 66.875 151.320 ;
        RECT 64.435 150.790 64.605 150.960 ;
        RECT 65.570 150.830 65.740 151.000 ;
        RECT 64.435 150.430 64.605 150.600 ;
        RECT 66.705 150.790 66.875 150.960 ;
        RECT 64.435 150.070 64.605 150.240 ;
        RECT 66.155 150.410 66.325 150.580 ;
        RECT 65.570 150.050 65.740 150.220 ;
        RECT 66.155 150.050 66.325 150.220 ;
        RECT 64.435 149.710 64.605 149.880 ;
        RECT 66.155 149.690 66.325 149.860 ;
        RECT 66.705 150.430 66.875 150.600 ;
        RECT 66.705 150.070 66.875 150.240 ;
        RECT 66.705 149.710 66.875 149.880 ;
        RECT 64.435 149.350 64.605 149.520 ;
        RECT 65.570 149.270 65.740 149.440 ;
        RECT 66.705 149.350 66.875 149.520 ;
        RECT 64.435 148.990 64.605 149.160 ;
        RECT 64.435 148.630 64.605 148.800 ;
        RECT 64.435 148.270 64.605 148.440 ;
        RECT 64.435 147.910 64.605 148.080 ;
        RECT 64.435 147.550 64.605 147.720 ;
        RECT 64.985 148.850 65.155 149.020 ;
        RECT 64.985 148.490 65.155 148.660 ;
        RECT 64.985 148.130 65.155 148.300 ;
        RECT 64.985 147.770 65.155 147.940 ;
        RECT 64.985 147.410 65.155 147.580 ;
        RECT 66.705 148.990 66.875 149.160 ;
        RECT 66.705 148.630 66.875 148.800 ;
        RECT 66.705 148.270 66.875 148.440 ;
        RECT 66.705 147.910 66.875 148.080 ;
        RECT 66.705 147.550 66.875 147.720 ;
        RECT 64.435 147.190 64.605 147.360 ;
        RECT 66.705 147.190 66.875 147.360 ;
        RECT 64.435 146.830 64.605 147.000 ;
        RECT 65.570 146.990 65.740 147.160 ;
        RECT 66.705 146.830 66.875 147.000 ;
        RECT 64.435 146.470 64.605 146.640 ;
        RECT 64.435 146.110 64.605 146.280 ;
        RECT 64.435 145.750 64.605 145.920 ;
        RECT 64.435 145.390 64.605 145.560 ;
        RECT 64.435 145.030 64.605 145.200 ;
        RECT 64.985 146.570 65.155 146.740 ;
        RECT 64.985 146.210 65.155 146.380 ;
        RECT 64.985 145.850 65.155 146.020 ;
        RECT 64.985 145.490 65.155 145.660 ;
        RECT 64.985 145.130 65.155 145.300 ;
        RECT 66.705 146.470 66.875 146.640 ;
        RECT 66.705 146.110 66.875 146.280 ;
        RECT 66.705 145.750 66.875 145.920 ;
        RECT 66.705 145.390 66.875 145.560 ;
        RECT 66.705 145.030 66.875 145.200 ;
        RECT 64.435 144.670 64.605 144.840 ;
        RECT 65.570 144.710 65.740 144.880 ;
        RECT 64.435 144.310 64.605 144.480 ;
        RECT 66.705 144.670 66.875 144.840 ;
        RECT 64.435 143.950 64.605 144.120 ;
        RECT 66.155 144.290 66.325 144.460 ;
        RECT 65.570 143.930 65.740 144.100 ;
        RECT 66.155 143.930 66.325 144.100 ;
        RECT 64.435 143.590 64.605 143.760 ;
        RECT 66.155 143.570 66.325 143.740 ;
        RECT 66.705 144.310 66.875 144.480 ;
        RECT 66.705 143.950 66.875 144.120 ;
        RECT 66.705 143.590 66.875 143.760 ;
        RECT 64.435 143.230 64.605 143.400 ;
        RECT 65.570 143.150 65.740 143.320 ;
        RECT 66.705 143.230 66.875 143.400 ;
        RECT 64.435 142.870 64.605 143.040 ;
        RECT 66.705 142.870 66.875 143.040 ;
        RECT 92.215 151.500 92.385 151.670 ;
        RECT 92.575 151.500 92.745 151.670 ;
        RECT 92.935 151.500 93.105 151.670 ;
        RECT 93.295 151.500 93.465 151.670 ;
        RECT 93.655 151.500 93.825 151.670 ;
        RECT 91.915 151.150 92.085 151.320 ;
        RECT 94.185 151.150 94.355 151.320 ;
        RECT 91.915 150.790 92.085 150.960 ;
        RECT 93.050 150.830 93.220 151.000 ;
        RECT 91.915 150.430 92.085 150.600 ;
        RECT 94.185 150.790 94.355 150.960 ;
        RECT 91.915 150.070 92.085 150.240 ;
        RECT 91.915 149.710 92.085 149.880 ;
        RECT 92.465 150.410 92.635 150.580 ;
        RECT 94.185 150.430 94.355 150.600 ;
        RECT 92.465 150.050 92.635 150.220 ;
        RECT 93.050 150.050 93.220 150.220 ;
        RECT 94.185 150.070 94.355 150.240 ;
        RECT 92.465 149.690 92.635 149.860 ;
        RECT 94.185 149.710 94.355 149.880 ;
        RECT 91.915 149.350 92.085 149.520 ;
        RECT 93.050 149.270 93.220 149.440 ;
        RECT 94.185 149.350 94.355 149.520 ;
        RECT 91.915 148.990 92.085 149.160 ;
        RECT 91.915 148.630 92.085 148.800 ;
        RECT 91.915 148.270 92.085 148.440 ;
        RECT 91.915 147.910 92.085 148.080 ;
        RECT 91.915 147.550 92.085 147.720 ;
        RECT 93.635 148.850 93.805 149.020 ;
        RECT 93.635 148.490 93.805 148.660 ;
        RECT 93.635 148.130 93.805 148.300 ;
        RECT 93.635 147.770 93.805 147.940 ;
        RECT 93.635 147.410 93.805 147.580 ;
        RECT 94.185 148.990 94.355 149.160 ;
        RECT 94.185 148.630 94.355 148.800 ;
        RECT 94.185 148.270 94.355 148.440 ;
        RECT 94.185 147.910 94.355 148.080 ;
        RECT 94.185 147.550 94.355 147.720 ;
        RECT 91.915 147.190 92.085 147.360 ;
        RECT 94.185 147.190 94.355 147.360 ;
        RECT 91.915 146.830 92.085 147.000 ;
        RECT 93.050 146.990 93.220 147.160 ;
        RECT 94.185 146.830 94.355 147.000 ;
        RECT 91.915 146.470 92.085 146.640 ;
        RECT 91.915 146.110 92.085 146.280 ;
        RECT 91.915 145.750 92.085 145.920 ;
        RECT 91.915 145.390 92.085 145.560 ;
        RECT 91.915 145.030 92.085 145.200 ;
        RECT 93.635 146.570 93.805 146.740 ;
        RECT 93.635 146.210 93.805 146.380 ;
        RECT 93.635 145.850 93.805 146.020 ;
        RECT 93.635 145.490 93.805 145.660 ;
        RECT 93.635 145.130 93.805 145.300 ;
        RECT 94.185 146.470 94.355 146.640 ;
        RECT 94.185 146.110 94.355 146.280 ;
        RECT 94.185 145.750 94.355 145.920 ;
        RECT 94.185 145.390 94.355 145.560 ;
        RECT 94.185 145.030 94.355 145.200 ;
        RECT 91.915 144.670 92.085 144.840 ;
        RECT 93.050 144.710 93.220 144.880 ;
        RECT 91.915 144.310 92.085 144.480 ;
        RECT 94.185 144.670 94.355 144.840 ;
        RECT 91.915 143.950 92.085 144.120 ;
        RECT 91.915 143.590 92.085 143.760 ;
        RECT 92.465 144.290 92.635 144.460 ;
        RECT 94.185 144.310 94.355 144.480 ;
        RECT 92.465 143.930 92.635 144.100 ;
        RECT 93.050 143.930 93.220 144.100 ;
        RECT 94.185 143.950 94.355 144.120 ;
        RECT 92.465 143.570 92.635 143.740 ;
        RECT 94.185 143.590 94.355 143.760 ;
        RECT 91.915 143.230 92.085 143.400 ;
        RECT 93.050 143.150 93.220 143.320 ;
        RECT 94.185 143.230 94.355 143.400 ;
        RECT 64.965 142.480 65.135 142.650 ;
        RECT 65.325 142.480 65.495 142.650 ;
        RECT 65.685 142.480 65.855 142.650 ;
        RECT 66.045 142.480 66.215 142.650 ;
        RECT 66.405 142.480 66.575 142.650 ;
        RECT 72.980 142.780 73.150 142.950 ;
        RECT 73.340 142.780 73.510 142.950 ;
        RECT 73.700 142.780 73.870 142.950 ;
        RECT 74.060 142.780 74.230 142.950 ;
        RECT 74.420 142.780 74.590 142.950 ;
        RECT 74.780 142.780 74.950 142.950 ;
        RECT 75.140 142.780 75.310 142.950 ;
        RECT 75.500 142.780 75.670 142.950 ;
        RECT 75.860 142.780 76.030 142.950 ;
        RECT 76.220 142.780 76.390 142.950 ;
        RECT 76.580 142.780 76.750 142.950 ;
        RECT 76.940 142.780 77.110 142.950 ;
        RECT 77.300 142.780 77.470 142.950 ;
        RECT 62.540 142.150 62.710 142.320 ;
        RECT 56.180 141.790 56.350 141.960 ;
        RECT 62.540 141.790 62.710 141.960 ;
        RECT 56.180 141.430 56.350 141.600 ;
        RECT 57.385 141.590 57.555 141.760 ;
        RECT 57.745 141.590 57.915 141.760 ;
        RECT 60.975 141.590 61.145 141.760 ;
        RECT 61.335 141.590 61.505 141.760 ;
        RECT 62.540 141.430 62.710 141.600 ;
        RECT 56.180 141.070 56.350 141.240 ;
        RECT 56.180 140.710 56.350 140.880 ;
        RECT 56.180 140.350 56.350 140.520 ;
        RECT 56.180 139.990 56.350 140.160 ;
        RECT 56.180 139.630 56.350 139.800 ;
        RECT 58.400 141.170 58.570 141.340 ;
        RECT 58.400 140.810 58.570 140.980 ;
        RECT 58.400 140.450 58.570 140.620 ;
        RECT 58.400 140.090 58.570 140.260 ;
        RECT 58.400 139.730 58.570 139.900 ;
        RECT 60.320 141.170 60.490 141.340 ;
        RECT 60.320 140.810 60.490 140.980 ;
        RECT 60.320 140.450 60.490 140.620 ;
        RECT 60.320 140.090 60.490 140.260 ;
        RECT 60.320 139.730 60.490 139.900 ;
        RECT 61.990 141.170 62.160 141.340 ;
        RECT 61.990 140.810 62.160 140.980 ;
        RECT 61.990 140.450 62.160 140.620 ;
        RECT 61.990 140.090 62.160 140.260 ;
        RECT 61.990 139.730 62.160 139.900 ;
        RECT 62.540 141.070 62.710 141.240 ;
        RECT 62.540 140.710 62.710 140.880 ;
        RECT 62.540 140.350 62.710 140.520 ;
        RECT 62.540 139.990 62.710 140.160 ;
        RECT 62.540 139.630 62.710 139.800 ;
        RECT 56.180 139.270 56.350 139.440 ;
        RECT 57.385 139.310 57.555 139.480 ;
        RECT 57.745 139.310 57.915 139.480 ;
        RECT 60.975 139.310 61.145 139.480 ;
        RECT 61.335 139.310 61.505 139.480 ;
        RECT 56.180 138.910 56.350 139.080 ;
        RECT 62.540 139.270 62.710 139.440 ;
        RECT 56.180 138.550 56.350 138.720 ;
        RECT 56.180 138.190 56.350 138.360 ;
        RECT 56.180 137.830 56.350 138.000 ;
        RECT 56.180 137.470 56.350 137.640 ;
        RECT 58.400 138.890 58.570 139.060 ;
        RECT 58.400 138.530 58.570 138.700 ;
        RECT 58.400 138.170 58.570 138.340 ;
        RECT 58.400 137.810 58.570 137.980 ;
        RECT 58.400 137.450 58.570 137.620 ;
        RECT 60.320 138.890 60.490 139.060 ;
        RECT 60.320 138.530 60.490 138.700 ;
        RECT 60.320 138.170 60.490 138.340 ;
        RECT 60.320 137.810 60.490 137.980 ;
        RECT 60.320 137.450 60.490 137.620 ;
        RECT 61.990 138.890 62.160 139.060 ;
        RECT 61.990 138.530 62.160 138.700 ;
        RECT 61.990 138.170 62.160 138.340 ;
        RECT 61.990 137.810 62.160 137.980 ;
        RECT 61.990 137.450 62.160 137.620 ;
        RECT 62.540 138.910 62.710 139.080 ;
        RECT 62.540 138.550 62.710 138.720 ;
        RECT 72.590 142.430 72.760 142.600 ;
        RECT 77.600 142.430 77.770 142.600 ;
        RECT 72.590 142.070 72.760 142.240 ;
        RECT 73.725 142.150 73.895 142.320 ;
        RECT 77.600 142.070 77.770 142.240 ;
        RECT 72.590 141.710 72.760 141.880 ;
        RECT 72.590 141.350 72.760 141.520 ;
        RECT 72.590 140.990 72.760 141.160 ;
        RECT 74.310 141.765 74.480 141.935 ;
        RECT 76.465 141.750 76.635 141.920 ;
        RECT 74.310 141.405 74.480 141.575 ;
        RECT 77.600 141.710 77.770 141.880 ;
        RECT 74.310 141.045 74.480 141.215 ;
        RECT 73.725 140.870 73.895 141.040 ;
        RECT 72.590 140.630 72.760 140.800 ;
        RECT 72.590 140.270 72.760 140.440 ;
        RECT 72.590 139.910 72.760 140.080 ;
        RECT 74.310 140.685 74.480 140.855 ;
        RECT 74.310 140.325 74.480 140.495 ;
        RECT 74.310 139.965 74.480 140.135 ;
        RECT 75.880 141.365 76.050 141.535 ;
        RECT 75.880 141.005 76.050 141.175 ;
        RECT 75.880 140.645 76.050 140.815 ;
        RECT 75.880 140.285 76.050 140.455 ;
        RECT 75.880 139.925 76.050 140.095 ;
        RECT 72.590 139.550 72.760 139.720 ;
        RECT 73.725 139.590 73.895 139.760 ;
        RECT 72.590 139.190 72.760 139.360 ;
        RECT 75.880 139.565 76.050 139.735 ;
        RECT 72.590 138.830 72.760 139.000 ;
        RECT 72.590 138.470 72.760 138.640 ;
        RECT 62.540 138.190 62.710 138.360 ;
        RECT 62.540 137.830 62.710 138.000 ;
        RECT 62.540 137.470 62.710 137.640 ;
        RECT 56.180 137.110 56.350 137.280 ;
        RECT 57.385 137.030 57.555 137.200 ;
        RECT 57.745 137.030 57.915 137.200 ;
        RECT 60.975 137.030 61.145 137.200 ;
        RECT 61.335 137.030 61.505 137.200 ;
        RECT 62.540 137.110 62.710 137.280 ;
        RECT 56.180 136.750 56.350 136.920 ;
        RECT 56.180 136.390 56.350 136.560 ;
        RECT 56.180 136.030 56.350 136.200 ;
        RECT 56.180 135.670 56.350 135.840 ;
        RECT 56.180 135.310 56.350 135.480 ;
        RECT 58.400 136.610 58.570 136.780 ;
        RECT 58.400 136.250 58.570 136.420 ;
        RECT 58.400 135.890 58.570 136.060 ;
        RECT 58.400 135.530 58.570 135.700 ;
        RECT 58.400 135.170 58.570 135.340 ;
        RECT 60.320 136.610 60.490 136.780 ;
        RECT 60.320 136.250 60.490 136.420 ;
        RECT 60.320 135.890 60.490 136.060 ;
        RECT 60.320 135.530 60.490 135.700 ;
        RECT 60.320 135.170 60.490 135.340 ;
        RECT 61.990 136.610 62.160 136.780 ;
        RECT 61.990 136.250 62.160 136.420 ;
        RECT 61.990 135.890 62.160 136.060 ;
        RECT 61.990 135.530 62.160 135.700 ;
        RECT 61.990 135.170 62.160 135.340 ;
        RECT 62.540 136.750 62.710 136.920 ;
        RECT 62.540 136.390 62.710 136.560 ;
        RECT 62.540 136.030 62.710 136.200 ;
        RECT 62.540 135.670 62.710 135.840 ;
        RECT 62.540 135.310 62.710 135.480 ;
        RECT 56.180 134.950 56.350 135.120 ;
        RECT 62.540 134.950 62.710 135.120 ;
        RECT 56.180 134.590 56.350 134.760 ;
        RECT 57.385 134.750 57.555 134.920 ;
        RECT 57.745 134.750 57.915 134.920 ;
        RECT 60.975 134.750 61.145 134.920 ;
        RECT 61.335 134.750 61.505 134.920 ;
        RECT 62.540 134.590 62.710 134.760 ;
        RECT 56.180 134.230 56.350 134.400 ;
        RECT 56.180 133.870 56.350 134.040 ;
        RECT 56.180 133.510 56.350 133.680 ;
        RECT 56.180 133.150 56.350 133.320 ;
        RECT 56.180 132.790 56.350 132.960 ;
        RECT 58.400 134.330 58.570 134.500 ;
        RECT 58.400 133.970 58.570 134.140 ;
        RECT 58.400 133.610 58.570 133.780 ;
        RECT 58.400 133.250 58.570 133.420 ;
        RECT 58.400 132.890 58.570 133.060 ;
        RECT 60.320 134.330 60.490 134.500 ;
        RECT 60.320 133.970 60.490 134.140 ;
        RECT 60.320 133.610 60.490 133.780 ;
        RECT 60.320 133.250 60.490 133.420 ;
        RECT 60.320 132.890 60.490 133.060 ;
        RECT 61.990 134.330 62.160 134.500 ;
        RECT 61.990 133.970 62.160 134.140 ;
        RECT 61.990 133.610 62.160 133.780 ;
        RECT 61.990 133.250 62.160 133.420 ;
        RECT 61.990 132.890 62.160 133.060 ;
        RECT 62.540 134.230 62.710 134.400 ;
        RECT 62.540 133.870 62.710 134.040 ;
        RECT 62.540 133.510 62.710 133.680 ;
        RECT 62.540 133.150 62.710 133.320 ;
        RECT 62.540 132.790 62.710 132.960 ;
        RECT 56.180 132.430 56.350 132.600 ;
        RECT 57.385 132.470 57.555 132.640 ;
        RECT 57.745 132.470 57.915 132.640 ;
        RECT 60.975 132.470 61.145 132.640 ;
        RECT 61.335 132.470 61.505 132.640 ;
        RECT 56.180 132.070 56.350 132.240 ;
        RECT 62.540 132.430 62.710 132.600 ;
        RECT 56.180 131.710 56.350 131.880 ;
        RECT 56.180 131.350 56.350 131.520 ;
        RECT 56.180 130.990 56.350 131.160 ;
        RECT 56.180 130.630 56.350 130.800 ;
        RECT 58.400 132.050 58.570 132.220 ;
        RECT 58.400 131.690 58.570 131.860 ;
        RECT 58.400 131.330 58.570 131.500 ;
        RECT 58.400 130.970 58.570 131.140 ;
        RECT 58.400 130.610 58.570 130.780 ;
        RECT 60.320 132.050 60.490 132.220 ;
        RECT 60.320 131.690 60.490 131.860 ;
        RECT 60.320 131.330 60.490 131.500 ;
        RECT 60.320 130.970 60.490 131.140 ;
        RECT 60.320 130.610 60.490 130.780 ;
        RECT 61.990 132.050 62.160 132.220 ;
        RECT 61.990 131.690 62.160 131.860 ;
        RECT 61.990 131.330 62.160 131.500 ;
        RECT 61.990 130.970 62.160 131.140 ;
        RECT 61.990 130.610 62.160 130.780 ;
        RECT 62.540 132.070 62.710 132.240 ;
        RECT 62.540 131.710 62.710 131.880 ;
        RECT 62.540 131.350 62.710 131.520 ;
        RECT 62.540 130.990 62.710 131.160 ;
        RECT 62.540 130.630 62.710 130.800 ;
        RECT 56.180 130.270 56.350 130.440 ;
        RECT 57.385 130.190 57.555 130.360 ;
        RECT 57.745 130.190 57.915 130.360 ;
        RECT 60.975 130.190 61.145 130.360 ;
        RECT 61.335 130.190 61.505 130.360 ;
        RECT 62.540 130.270 62.710 130.440 ;
        RECT 56.180 129.910 56.350 130.080 ;
        RECT 56.180 129.550 56.350 129.720 ;
        RECT 56.180 129.190 56.350 129.360 ;
        RECT 56.180 128.830 56.350 129.000 ;
        RECT 56.180 128.470 56.350 128.640 ;
        RECT 56.730 129.770 56.900 129.940 ;
        RECT 56.730 129.410 56.900 129.580 ;
        RECT 56.730 129.050 56.900 129.220 ;
        RECT 56.730 128.690 56.900 128.860 ;
        RECT 56.730 128.330 56.900 128.500 ;
        RECT 60.320 129.770 60.490 129.940 ;
        RECT 60.320 129.410 60.490 129.580 ;
        RECT 60.320 129.050 60.490 129.220 ;
        RECT 60.320 128.690 60.490 128.860 ;
        RECT 60.320 128.330 60.490 128.500 ;
        RECT 61.990 129.770 62.160 129.940 ;
        RECT 61.990 129.410 62.160 129.580 ;
        RECT 61.990 129.050 62.160 129.220 ;
        RECT 61.990 128.690 62.160 128.860 ;
        RECT 61.990 128.330 62.160 128.500 ;
        RECT 62.540 129.910 62.710 130.080 ;
        RECT 62.540 129.550 62.710 129.720 ;
        RECT 62.540 129.190 62.710 129.360 ;
        RECT 62.540 128.830 62.710 129.000 ;
        RECT 62.540 128.470 62.710 128.640 ;
        RECT 56.180 128.110 56.350 128.280 ;
        RECT 62.540 128.110 62.710 128.280 ;
        RECT 56.180 127.750 56.350 127.920 ;
        RECT 57.385 127.910 57.555 128.080 ;
        RECT 57.745 127.910 57.915 128.080 ;
        RECT 60.975 127.910 61.145 128.080 ;
        RECT 61.335 127.910 61.505 128.080 ;
        RECT 62.540 127.750 62.710 127.920 ;
        RECT 56.180 127.390 56.350 127.560 ;
        RECT 56.180 127.030 56.350 127.200 ;
        RECT 56.180 126.670 56.350 126.840 ;
        RECT 56.180 126.310 56.350 126.480 ;
        RECT 56.180 125.950 56.350 126.120 ;
        RECT 56.730 127.490 56.900 127.660 ;
        RECT 56.730 127.130 56.900 127.300 ;
        RECT 56.730 126.770 56.900 126.940 ;
        RECT 56.730 126.410 56.900 126.580 ;
        RECT 56.730 126.050 56.900 126.220 ;
        RECT 60.320 127.490 60.490 127.660 ;
        RECT 60.320 127.130 60.490 127.300 ;
        RECT 60.320 126.770 60.490 126.940 ;
        RECT 60.320 126.410 60.490 126.580 ;
        RECT 60.320 126.050 60.490 126.220 ;
        RECT 61.990 127.490 62.160 127.660 ;
        RECT 61.990 127.130 62.160 127.300 ;
        RECT 61.990 126.770 62.160 126.940 ;
        RECT 61.990 126.410 62.160 126.580 ;
        RECT 61.990 126.050 62.160 126.220 ;
        RECT 62.540 127.390 62.710 127.560 ;
        RECT 62.540 127.030 62.710 127.200 ;
        RECT 62.540 126.670 62.710 126.840 ;
        RECT 62.540 126.310 62.710 126.480 ;
        RECT 62.540 125.950 62.710 126.120 ;
        RECT 56.180 125.590 56.350 125.760 ;
        RECT 57.385 125.630 57.555 125.800 ;
        RECT 57.745 125.630 57.915 125.800 ;
        RECT 60.975 125.630 61.145 125.800 ;
        RECT 61.335 125.630 61.505 125.800 ;
        RECT 56.180 125.230 56.350 125.400 ;
        RECT 62.540 125.590 62.710 125.760 ;
        RECT 56.180 124.870 56.350 125.040 ;
        RECT 56.180 124.510 56.350 124.680 ;
        RECT 56.180 124.150 56.350 124.320 ;
        RECT 56.180 123.790 56.350 123.960 ;
        RECT 58.400 125.210 58.570 125.380 ;
        RECT 58.400 124.850 58.570 125.020 ;
        RECT 58.400 124.490 58.570 124.660 ;
        RECT 58.400 124.130 58.570 124.300 ;
        RECT 58.400 123.770 58.570 123.940 ;
        RECT 60.320 125.210 60.490 125.380 ;
        RECT 60.320 124.850 60.490 125.020 ;
        RECT 60.320 124.490 60.490 124.660 ;
        RECT 60.320 124.130 60.490 124.300 ;
        RECT 60.320 123.770 60.490 123.940 ;
        RECT 61.990 125.210 62.160 125.380 ;
        RECT 61.990 124.850 62.160 125.020 ;
        RECT 61.990 124.490 62.160 124.660 ;
        RECT 61.990 124.130 62.160 124.300 ;
        RECT 61.990 123.770 62.160 123.940 ;
        RECT 62.540 125.230 62.710 125.400 ;
        RECT 62.540 124.870 62.710 125.040 ;
        RECT 62.540 124.510 62.710 124.680 ;
        RECT 62.540 124.150 62.710 124.320 ;
        RECT 62.540 123.790 62.710 123.960 ;
        RECT 56.180 123.430 56.350 123.600 ;
        RECT 57.385 123.350 57.555 123.520 ;
        RECT 57.745 123.350 57.915 123.520 ;
        RECT 60.975 123.350 61.145 123.520 ;
        RECT 61.335 123.350 61.505 123.520 ;
        RECT 62.540 123.430 62.710 123.600 ;
        RECT 56.180 123.070 56.350 123.240 ;
        RECT 56.180 122.710 56.350 122.880 ;
        RECT 56.180 122.350 56.350 122.520 ;
        RECT 56.180 121.990 56.350 122.160 ;
        RECT 56.180 121.630 56.350 121.800 ;
        RECT 58.400 122.930 58.570 123.100 ;
        RECT 58.400 122.570 58.570 122.740 ;
        RECT 58.400 122.210 58.570 122.380 ;
        RECT 58.400 121.850 58.570 122.020 ;
        RECT 58.400 121.490 58.570 121.660 ;
        RECT 60.320 122.930 60.490 123.100 ;
        RECT 60.320 122.570 60.490 122.740 ;
        RECT 60.320 122.210 60.490 122.380 ;
        RECT 60.320 121.850 60.490 122.020 ;
        RECT 60.320 121.490 60.490 121.660 ;
        RECT 61.990 122.930 62.160 123.100 ;
        RECT 61.990 122.570 62.160 122.740 ;
        RECT 61.990 122.210 62.160 122.380 ;
        RECT 61.990 121.850 62.160 122.020 ;
        RECT 61.990 121.490 62.160 121.660 ;
        RECT 62.540 123.070 62.710 123.240 ;
        RECT 62.540 122.710 62.710 122.880 ;
        RECT 62.540 122.350 62.710 122.520 ;
        RECT 62.540 121.990 62.710 122.160 ;
        RECT 62.540 121.630 62.710 121.800 ;
        RECT 56.180 121.270 56.350 121.440 ;
        RECT 62.540 121.270 62.710 121.440 ;
        RECT 56.180 120.910 56.350 121.080 ;
        RECT 57.385 121.070 57.555 121.240 ;
        RECT 57.745 121.070 57.915 121.240 ;
        RECT 60.975 121.070 61.145 121.240 ;
        RECT 61.335 121.070 61.505 121.240 ;
        RECT 62.540 120.910 62.710 121.080 ;
        RECT 56.180 120.550 56.350 120.720 ;
        RECT 56.180 120.190 56.350 120.360 ;
        RECT 56.180 119.830 56.350 120.000 ;
        RECT 56.180 119.470 56.350 119.640 ;
        RECT 56.180 119.110 56.350 119.280 ;
        RECT 58.400 120.650 58.570 120.820 ;
        RECT 58.400 120.290 58.570 120.460 ;
        RECT 58.400 119.930 58.570 120.100 ;
        RECT 58.400 119.570 58.570 119.740 ;
        RECT 58.400 119.210 58.570 119.380 ;
        RECT 60.320 120.650 60.490 120.820 ;
        RECT 60.320 120.290 60.490 120.460 ;
        RECT 60.320 119.930 60.490 120.100 ;
        RECT 60.320 119.570 60.490 119.740 ;
        RECT 60.320 119.210 60.490 119.380 ;
        RECT 61.990 120.650 62.160 120.820 ;
        RECT 61.990 120.290 62.160 120.460 ;
        RECT 61.990 119.930 62.160 120.100 ;
        RECT 61.990 119.570 62.160 119.740 ;
        RECT 61.990 119.210 62.160 119.380 ;
        RECT 62.540 120.550 62.710 120.720 ;
        RECT 62.540 120.190 62.710 120.360 ;
        RECT 62.540 119.830 62.710 120.000 ;
        RECT 62.540 119.470 62.710 119.640 ;
        RECT 62.540 119.110 62.710 119.280 ;
        RECT 56.180 118.750 56.350 118.920 ;
        RECT 57.385 118.790 57.555 118.960 ;
        RECT 57.745 118.790 57.915 118.960 ;
        RECT 60.975 118.790 61.145 118.960 ;
        RECT 61.335 118.790 61.505 118.960 ;
        RECT 56.180 118.390 56.350 118.560 ;
        RECT 62.540 118.750 62.710 118.920 ;
        RECT 56.180 118.030 56.350 118.200 ;
        RECT 56.180 117.670 56.350 117.840 ;
        RECT 56.180 117.310 56.350 117.480 ;
        RECT 56.180 116.950 56.350 117.120 ;
        RECT 58.400 118.370 58.570 118.540 ;
        RECT 58.400 118.010 58.570 118.180 ;
        RECT 58.400 117.650 58.570 117.820 ;
        RECT 58.400 117.290 58.570 117.460 ;
        RECT 58.400 116.930 58.570 117.100 ;
        RECT 60.320 118.370 60.490 118.540 ;
        RECT 60.320 118.010 60.490 118.180 ;
        RECT 60.320 117.650 60.490 117.820 ;
        RECT 60.320 117.290 60.490 117.460 ;
        RECT 60.320 116.930 60.490 117.100 ;
        RECT 61.990 118.370 62.160 118.540 ;
        RECT 61.990 118.010 62.160 118.180 ;
        RECT 61.990 117.650 62.160 117.820 ;
        RECT 61.990 117.290 62.160 117.460 ;
        RECT 61.990 116.930 62.160 117.100 ;
        RECT 62.540 118.390 62.710 118.560 ;
        RECT 62.540 118.030 62.710 118.200 ;
        RECT 62.540 117.670 62.710 117.840 ;
        RECT 64.965 138.290 65.135 138.460 ;
        RECT 65.325 138.290 65.495 138.460 ;
        RECT 65.685 138.290 65.855 138.460 ;
        RECT 66.045 138.290 66.215 138.460 ;
        RECT 66.405 138.290 66.575 138.460 ;
        RECT 64.435 137.940 64.605 138.110 ;
        RECT 66.705 137.940 66.875 138.110 ;
        RECT 64.435 137.580 64.605 137.750 ;
        RECT 65.570 137.620 65.740 137.790 ;
        RECT 66.705 137.580 66.875 137.750 ;
        RECT 64.435 137.220 64.605 137.390 ;
        RECT 64.435 136.860 64.605 137.030 ;
        RECT 64.435 136.500 64.605 136.670 ;
        RECT 64.435 136.140 64.605 136.310 ;
        RECT 64.435 135.780 64.605 135.950 ;
        RECT 64.435 135.420 64.605 135.590 ;
        RECT 64.985 137.235 65.155 137.405 ;
        RECT 64.985 136.875 65.155 137.045 ;
        RECT 64.985 136.515 65.155 136.685 ;
        RECT 66.155 137.235 66.325 137.405 ;
        RECT 66.155 136.875 66.325 137.045 ;
        RECT 66.155 136.515 66.325 136.685 ;
        RECT 65.570 136.340 65.740 136.510 ;
        RECT 64.985 136.155 65.155 136.325 ;
        RECT 64.985 135.795 65.155 135.965 ;
        RECT 64.985 135.435 65.155 135.605 ;
        RECT 66.155 136.155 66.325 136.325 ;
        RECT 66.155 135.795 66.325 135.965 ;
        RECT 66.155 135.435 66.325 135.605 ;
        RECT 66.705 137.220 66.875 137.390 ;
        RECT 66.705 136.860 66.875 137.030 ;
        RECT 66.705 136.500 66.875 136.670 ;
        RECT 66.705 136.140 66.875 136.310 ;
        RECT 66.705 135.780 66.875 135.950 ;
        RECT 66.705 135.420 66.875 135.590 ;
        RECT 64.435 135.060 64.605 135.230 ;
        RECT 65.570 135.060 65.740 135.230 ;
        RECT 66.705 135.060 66.875 135.230 ;
        RECT 64.435 134.700 64.605 134.870 ;
        RECT 64.435 134.340 64.605 134.510 ;
        RECT 64.435 133.980 64.605 134.150 ;
        RECT 64.435 133.620 64.605 133.790 ;
        RECT 64.435 133.260 64.605 133.430 ;
        RECT 64.985 134.640 65.155 134.810 ;
        RECT 64.985 134.280 65.155 134.450 ;
        RECT 64.985 133.920 65.155 134.090 ;
        RECT 64.985 133.560 65.155 133.730 ;
        RECT 64.985 133.200 65.155 133.370 ;
        RECT 66.155 134.640 66.325 134.810 ;
        RECT 66.155 134.280 66.325 134.450 ;
        RECT 66.155 133.920 66.325 134.090 ;
        RECT 66.155 133.560 66.325 133.730 ;
        RECT 66.155 133.200 66.325 133.370 ;
        RECT 66.705 134.700 66.875 134.870 ;
        RECT 66.705 134.340 66.875 134.510 ;
        RECT 66.705 133.980 66.875 134.150 ;
        RECT 66.705 133.620 66.875 133.790 ;
        RECT 66.705 133.260 66.875 133.430 ;
        RECT 64.435 132.900 64.605 133.070 ;
        RECT 65.570 132.780 65.740 132.950 ;
        RECT 66.705 132.900 66.875 133.070 ;
        RECT 64.435 132.540 64.605 132.710 ;
        RECT 66.705 132.540 66.875 132.710 ;
        RECT 64.435 132.180 64.605 132.350 ;
        RECT 64.435 131.820 64.605 131.990 ;
        RECT 64.435 131.460 64.605 131.630 ;
        RECT 64.435 131.100 64.605 131.270 ;
        RECT 64.985 132.360 65.155 132.530 ;
        RECT 64.985 132.000 65.155 132.170 ;
        RECT 64.985 131.640 65.155 131.810 ;
        RECT 64.985 131.280 65.155 131.450 ;
        RECT 64.985 130.920 65.155 131.090 ;
        RECT 66.155 132.360 66.325 132.530 ;
        RECT 66.155 132.000 66.325 132.170 ;
        RECT 66.155 131.640 66.325 131.810 ;
        RECT 66.155 131.280 66.325 131.450 ;
        RECT 66.155 130.920 66.325 131.090 ;
        RECT 66.705 132.180 66.875 132.350 ;
        RECT 66.705 131.820 66.875 131.990 ;
        RECT 66.705 131.460 66.875 131.630 ;
        RECT 66.705 131.100 66.875 131.270 ;
        RECT 64.435 130.740 64.605 130.910 ;
        RECT 66.705 130.740 66.875 130.910 ;
        RECT 64.435 130.380 64.605 130.550 ;
        RECT 65.570 130.500 65.740 130.670 ;
        RECT 66.705 130.380 66.875 130.550 ;
        RECT 64.435 130.020 64.605 130.190 ;
        RECT 64.435 129.660 64.605 129.830 ;
        RECT 64.435 129.300 64.605 129.470 ;
        RECT 64.435 128.940 64.605 129.110 ;
        RECT 64.435 128.580 64.605 128.750 ;
        RECT 64.435 128.220 64.605 128.390 ;
        RECT 64.985 130.115 65.155 130.285 ;
        RECT 64.985 129.755 65.155 129.925 ;
        RECT 64.985 129.395 65.155 129.565 ;
        RECT 66.155 130.115 66.325 130.285 ;
        RECT 66.155 129.755 66.325 129.925 ;
        RECT 66.155 129.395 66.325 129.565 ;
        RECT 65.570 129.220 65.740 129.390 ;
        RECT 64.985 129.035 65.155 129.205 ;
        RECT 64.985 128.675 65.155 128.845 ;
        RECT 64.985 128.315 65.155 128.485 ;
        RECT 66.155 129.035 66.325 129.205 ;
        RECT 66.155 128.675 66.325 128.845 ;
        RECT 66.155 128.315 66.325 128.485 ;
        RECT 66.705 130.020 66.875 130.190 ;
        RECT 66.705 129.660 66.875 129.830 ;
        RECT 66.705 129.300 66.875 129.470 ;
        RECT 66.705 128.940 66.875 129.110 ;
        RECT 66.705 128.580 66.875 128.750 ;
        RECT 66.705 128.220 66.875 128.390 ;
        RECT 64.435 127.860 64.605 128.030 ;
        RECT 65.570 127.940 65.740 128.110 ;
        RECT 66.705 127.860 66.875 128.030 ;
        RECT 64.435 127.500 64.605 127.670 ;
        RECT 64.435 127.140 64.605 127.310 ;
        RECT 64.435 126.780 64.605 126.950 ;
        RECT 64.435 126.420 64.605 126.590 ;
        RECT 64.435 126.060 64.605 126.230 ;
        RECT 64.435 125.700 64.605 125.870 ;
        RECT 64.985 127.555 65.155 127.725 ;
        RECT 64.985 127.195 65.155 127.365 ;
        RECT 64.985 126.835 65.155 127.005 ;
        RECT 66.155 127.555 66.325 127.725 ;
        RECT 66.155 127.195 66.325 127.365 ;
        RECT 66.155 126.835 66.325 127.005 ;
        RECT 65.570 126.660 65.740 126.830 ;
        RECT 64.985 126.475 65.155 126.645 ;
        RECT 64.985 126.115 65.155 126.285 ;
        RECT 64.985 125.755 65.155 125.925 ;
        RECT 66.155 126.475 66.325 126.645 ;
        RECT 66.155 126.115 66.325 126.285 ;
        RECT 66.155 125.755 66.325 125.925 ;
        RECT 66.705 127.500 66.875 127.670 ;
        RECT 66.705 127.140 66.875 127.310 ;
        RECT 66.705 126.780 66.875 126.950 ;
        RECT 66.705 126.420 66.875 126.590 ;
        RECT 66.705 126.060 66.875 126.230 ;
        RECT 66.705 125.700 66.875 125.870 ;
        RECT 64.435 125.340 64.605 125.510 ;
        RECT 65.570 125.380 65.740 125.550 ;
        RECT 64.435 124.980 64.605 125.150 ;
        RECT 66.705 125.340 66.875 125.510 ;
        RECT 64.435 124.620 64.605 124.790 ;
        RECT 64.435 124.260 64.605 124.430 ;
        RECT 64.435 123.900 64.605 124.070 ;
        RECT 64.435 123.540 64.605 123.710 ;
        RECT 64.985 124.960 65.155 125.130 ;
        RECT 64.985 124.600 65.155 124.770 ;
        RECT 64.985 124.240 65.155 124.410 ;
        RECT 64.985 123.880 65.155 124.050 ;
        RECT 64.985 123.520 65.155 123.690 ;
        RECT 66.705 124.980 66.875 125.150 ;
        RECT 66.705 124.620 66.875 124.790 ;
        RECT 66.705 124.260 66.875 124.430 ;
        RECT 66.705 123.900 66.875 124.070 ;
        RECT 66.705 123.540 66.875 123.710 ;
        RECT 64.435 123.180 64.605 123.350 ;
        RECT 65.570 123.100 65.740 123.270 ;
        RECT 66.705 123.180 66.875 123.350 ;
        RECT 64.435 122.820 64.605 122.990 ;
        RECT 64.435 122.460 64.605 122.630 ;
        RECT 64.435 122.100 64.605 122.270 ;
        RECT 64.435 121.740 64.605 121.910 ;
        RECT 64.435 121.380 64.605 121.550 ;
        RECT 64.985 122.680 65.155 122.850 ;
        RECT 64.985 122.320 65.155 122.490 ;
        RECT 64.985 121.960 65.155 122.130 ;
        RECT 64.985 121.600 65.155 121.770 ;
        RECT 64.985 121.240 65.155 121.410 ;
        RECT 66.705 122.820 66.875 122.990 ;
        RECT 66.705 122.460 66.875 122.630 ;
        RECT 66.705 122.100 66.875 122.270 ;
        RECT 66.705 121.740 66.875 121.910 ;
        RECT 66.705 121.380 66.875 121.550 ;
        RECT 64.435 121.020 64.605 121.190 ;
        RECT 66.705 121.020 66.875 121.190 ;
        RECT 64.435 120.660 64.605 120.830 ;
        RECT 65.570 120.820 65.740 120.990 ;
        RECT 66.705 120.660 66.875 120.830 ;
        RECT 64.435 120.300 64.605 120.470 ;
        RECT 64.435 119.940 64.605 120.110 ;
        RECT 64.435 119.580 64.605 119.750 ;
        RECT 64.435 119.220 64.605 119.390 ;
        RECT 64.435 118.860 64.605 119.030 ;
        RECT 64.435 118.500 64.605 118.670 ;
        RECT 64.985 120.435 65.155 120.605 ;
        RECT 64.985 120.075 65.155 120.245 ;
        RECT 64.985 119.715 65.155 119.885 ;
        RECT 66.155 120.435 66.325 120.605 ;
        RECT 66.155 120.075 66.325 120.245 ;
        RECT 66.155 119.715 66.325 119.885 ;
        RECT 65.570 119.540 65.740 119.710 ;
        RECT 64.985 119.355 65.155 119.525 ;
        RECT 64.985 118.995 65.155 119.165 ;
        RECT 64.985 118.635 65.155 118.805 ;
        RECT 66.155 119.355 66.325 119.525 ;
        RECT 66.155 118.995 66.325 119.165 ;
        RECT 66.155 118.635 66.325 118.805 ;
        RECT 66.705 120.300 66.875 120.470 ;
        RECT 66.705 119.940 66.875 120.110 ;
        RECT 66.705 119.580 66.875 119.750 ;
        RECT 66.705 119.220 66.875 119.390 ;
        RECT 66.705 118.860 66.875 119.030 ;
        RECT 66.705 118.500 66.875 118.670 ;
        RECT 64.435 118.140 64.605 118.310 ;
        RECT 65.570 118.260 65.740 118.430 ;
        RECT 66.705 118.140 66.875 118.310 ;
        RECT 64.965 117.590 65.135 117.760 ;
        RECT 65.325 117.590 65.495 117.760 ;
        RECT 65.685 117.590 65.855 117.760 ;
        RECT 66.045 117.590 66.215 117.760 ;
        RECT 66.405 117.590 66.575 117.760 ;
        RECT 68.500 138.290 68.670 138.460 ;
        RECT 68.860 138.290 69.030 138.460 ;
        RECT 69.220 138.290 69.390 138.460 ;
        RECT 69.580 138.290 69.750 138.460 ;
        RECT 69.940 138.290 70.110 138.460 ;
        RECT 70.300 138.290 70.470 138.460 ;
        RECT 70.660 138.290 70.830 138.460 ;
        RECT 68.190 137.940 68.360 138.110 ;
        RECT 70.960 137.940 71.130 138.110 ;
        RECT 68.190 137.580 68.360 137.750 ;
        RECT 69.395 137.620 69.565 137.790 ;
        RECT 69.755 137.620 69.925 137.790 ;
        RECT 70.960 137.580 71.130 137.750 ;
        RECT 68.190 137.220 68.360 137.390 ;
        RECT 68.190 136.860 68.360 137.030 ;
        RECT 68.190 136.500 68.360 136.670 ;
        RECT 68.190 136.140 68.360 136.310 ;
        RECT 68.190 135.780 68.360 135.950 ;
        RECT 68.190 135.420 68.360 135.590 ;
        RECT 68.740 137.235 68.910 137.405 ;
        RECT 68.740 136.875 68.910 137.045 ;
        RECT 68.740 136.515 68.910 136.685 ;
        RECT 70.410 137.235 70.580 137.405 ;
        RECT 70.410 136.875 70.580 137.045 ;
        RECT 70.410 136.515 70.580 136.685 ;
        RECT 69.395 136.340 69.565 136.510 ;
        RECT 69.755 136.340 69.925 136.510 ;
        RECT 68.740 136.155 68.910 136.325 ;
        RECT 68.740 135.795 68.910 135.965 ;
        RECT 68.740 135.435 68.910 135.605 ;
        RECT 70.410 136.155 70.580 136.325 ;
        RECT 70.410 135.795 70.580 135.965 ;
        RECT 70.410 135.435 70.580 135.605 ;
        RECT 70.960 137.220 71.130 137.390 ;
        RECT 70.960 136.860 71.130 137.030 ;
        RECT 70.960 136.500 71.130 136.670 ;
        RECT 70.960 136.140 71.130 136.310 ;
        RECT 70.960 135.780 71.130 135.950 ;
        RECT 70.960 135.420 71.130 135.590 ;
        RECT 68.190 135.060 68.360 135.230 ;
        RECT 69.395 135.060 69.565 135.230 ;
        RECT 69.755 135.060 69.925 135.230 ;
        RECT 70.960 135.060 71.130 135.230 ;
        RECT 68.190 134.700 68.360 134.870 ;
        RECT 68.190 134.340 68.360 134.510 ;
        RECT 68.190 133.980 68.360 134.150 ;
        RECT 68.190 133.620 68.360 133.790 ;
        RECT 68.190 133.260 68.360 133.430 ;
        RECT 68.740 134.640 68.910 134.810 ;
        RECT 68.740 134.280 68.910 134.450 ;
        RECT 68.740 133.920 68.910 134.090 ;
        RECT 68.740 133.560 68.910 133.730 ;
        RECT 68.740 133.200 68.910 133.370 ;
        RECT 70.410 134.640 70.580 134.810 ;
        RECT 70.410 134.280 70.580 134.450 ;
        RECT 70.410 133.920 70.580 134.090 ;
        RECT 70.410 133.560 70.580 133.730 ;
        RECT 70.410 133.200 70.580 133.370 ;
        RECT 70.960 134.700 71.130 134.870 ;
        RECT 70.960 134.340 71.130 134.510 ;
        RECT 70.960 133.980 71.130 134.150 ;
        RECT 70.960 133.620 71.130 133.790 ;
        RECT 70.960 133.260 71.130 133.430 ;
        RECT 68.190 132.900 68.360 133.070 ;
        RECT 69.395 132.780 69.565 132.950 ;
        RECT 69.755 132.780 69.925 132.950 ;
        RECT 70.960 132.900 71.130 133.070 ;
        RECT 68.190 132.540 68.360 132.710 ;
        RECT 70.960 132.540 71.130 132.710 ;
        RECT 68.190 132.180 68.360 132.350 ;
        RECT 68.190 131.820 68.360 131.990 ;
        RECT 68.190 131.460 68.360 131.630 ;
        RECT 68.190 131.100 68.360 131.270 ;
        RECT 68.740 132.360 68.910 132.530 ;
        RECT 68.740 132.000 68.910 132.170 ;
        RECT 68.740 131.640 68.910 131.810 ;
        RECT 68.740 131.280 68.910 131.450 ;
        RECT 68.740 130.920 68.910 131.090 ;
        RECT 70.410 132.360 70.580 132.530 ;
        RECT 70.410 132.000 70.580 132.170 ;
        RECT 70.410 131.640 70.580 131.810 ;
        RECT 70.410 131.280 70.580 131.450 ;
        RECT 70.410 130.920 70.580 131.090 ;
        RECT 70.960 132.180 71.130 132.350 ;
        RECT 70.960 131.820 71.130 131.990 ;
        RECT 70.960 131.460 71.130 131.630 ;
        RECT 70.960 131.100 71.130 131.270 ;
        RECT 68.190 130.740 68.360 130.910 ;
        RECT 70.960 130.740 71.130 130.910 ;
        RECT 68.190 130.380 68.360 130.550 ;
        RECT 69.395 130.500 69.565 130.670 ;
        RECT 69.755 130.500 69.925 130.670 ;
        RECT 70.960 130.380 71.130 130.550 ;
        RECT 68.190 130.020 68.360 130.190 ;
        RECT 68.190 129.660 68.360 129.830 ;
        RECT 68.190 129.300 68.360 129.470 ;
        RECT 68.190 128.940 68.360 129.110 ;
        RECT 68.190 128.580 68.360 128.750 ;
        RECT 68.190 128.220 68.360 128.390 ;
        RECT 68.740 130.115 68.910 130.285 ;
        RECT 68.740 129.755 68.910 129.925 ;
        RECT 68.740 129.395 68.910 129.565 ;
        RECT 70.410 130.115 70.580 130.285 ;
        RECT 70.410 129.755 70.580 129.925 ;
        RECT 70.410 129.395 70.580 129.565 ;
        RECT 69.395 129.220 69.565 129.390 ;
        RECT 69.755 129.220 69.925 129.390 ;
        RECT 68.740 129.035 68.910 129.205 ;
        RECT 68.740 128.675 68.910 128.845 ;
        RECT 68.740 128.315 68.910 128.485 ;
        RECT 70.410 129.035 70.580 129.205 ;
        RECT 70.410 128.675 70.580 128.845 ;
        RECT 70.410 128.315 70.580 128.485 ;
        RECT 70.960 130.020 71.130 130.190 ;
        RECT 70.960 129.660 71.130 129.830 ;
        RECT 70.960 129.300 71.130 129.470 ;
        RECT 70.960 128.940 71.130 129.110 ;
        RECT 70.960 128.580 71.130 128.750 ;
        RECT 70.960 128.220 71.130 128.390 ;
        RECT 68.190 127.860 68.360 128.030 ;
        RECT 69.395 127.940 69.565 128.110 ;
        RECT 69.755 127.940 69.925 128.110 ;
        RECT 70.960 127.860 71.130 128.030 ;
        RECT 68.190 127.500 68.360 127.670 ;
        RECT 68.190 127.140 68.360 127.310 ;
        RECT 68.190 126.780 68.360 126.950 ;
        RECT 68.190 126.420 68.360 126.590 ;
        RECT 68.190 126.060 68.360 126.230 ;
        RECT 68.190 125.700 68.360 125.870 ;
        RECT 68.740 127.555 68.910 127.725 ;
        RECT 68.740 127.195 68.910 127.365 ;
        RECT 68.740 126.835 68.910 127.005 ;
        RECT 70.410 127.555 70.580 127.725 ;
        RECT 70.410 127.195 70.580 127.365 ;
        RECT 70.410 126.835 70.580 127.005 ;
        RECT 69.395 126.660 69.565 126.830 ;
        RECT 69.755 126.660 69.925 126.830 ;
        RECT 68.740 126.475 68.910 126.645 ;
        RECT 68.740 126.115 68.910 126.285 ;
        RECT 68.740 125.755 68.910 125.925 ;
        RECT 70.410 126.475 70.580 126.645 ;
        RECT 70.410 126.115 70.580 126.285 ;
        RECT 70.410 125.755 70.580 125.925 ;
        RECT 70.960 127.500 71.130 127.670 ;
        RECT 70.960 127.140 71.130 127.310 ;
        RECT 70.960 126.780 71.130 126.950 ;
        RECT 70.960 126.420 71.130 126.590 ;
        RECT 70.960 126.060 71.130 126.230 ;
        RECT 70.960 125.700 71.130 125.870 ;
        RECT 68.190 125.340 68.360 125.510 ;
        RECT 69.395 125.380 69.565 125.550 ;
        RECT 69.755 125.380 69.925 125.550 ;
        RECT 68.190 124.980 68.360 125.150 ;
        RECT 70.960 125.340 71.130 125.510 ;
        RECT 68.190 124.620 68.360 124.790 ;
        RECT 68.190 124.260 68.360 124.430 ;
        RECT 68.190 123.900 68.360 124.070 ;
        RECT 68.190 123.540 68.360 123.710 ;
        RECT 70.410 124.960 70.580 125.130 ;
        RECT 70.410 124.600 70.580 124.770 ;
        RECT 70.410 124.240 70.580 124.410 ;
        RECT 70.410 123.880 70.580 124.050 ;
        RECT 70.410 123.520 70.580 123.690 ;
        RECT 70.960 124.980 71.130 125.150 ;
        RECT 70.960 124.620 71.130 124.790 ;
        RECT 70.960 124.260 71.130 124.430 ;
        RECT 70.960 123.900 71.130 124.070 ;
        RECT 70.960 123.540 71.130 123.710 ;
        RECT 68.190 123.180 68.360 123.350 ;
        RECT 69.395 123.100 69.565 123.270 ;
        RECT 69.755 123.100 69.925 123.270 ;
        RECT 70.960 123.180 71.130 123.350 ;
        RECT 68.190 122.820 68.360 122.990 ;
        RECT 68.190 122.460 68.360 122.630 ;
        RECT 68.190 122.100 68.360 122.270 ;
        RECT 68.190 121.740 68.360 121.910 ;
        RECT 68.190 121.380 68.360 121.550 ;
        RECT 70.410 122.680 70.580 122.850 ;
        RECT 70.410 122.320 70.580 122.490 ;
        RECT 70.410 121.960 70.580 122.130 ;
        RECT 70.410 121.600 70.580 121.770 ;
        RECT 70.410 121.240 70.580 121.410 ;
        RECT 70.960 122.820 71.130 122.990 ;
        RECT 70.960 122.460 71.130 122.630 ;
        RECT 70.960 122.100 71.130 122.270 ;
        RECT 70.960 121.740 71.130 121.910 ;
        RECT 70.960 121.380 71.130 121.550 ;
        RECT 68.190 121.020 68.360 121.190 ;
        RECT 70.960 121.020 71.130 121.190 ;
        RECT 68.190 120.660 68.360 120.830 ;
        RECT 69.395 120.820 69.565 120.990 ;
        RECT 69.755 120.820 69.925 120.990 ;
        RECT 70.960 120.660 71.130 120.830 ;
        RECT 68.190 120.300 68.360 120.470 ;
        RECT 68.190 119.940 68.360 120.110 ;
        RECT 68.190 119.580 68.360 119.750 ;
        RECT 68.190 119.220 68.360 119.390 ;
        RECT 68.190 118.860 68.360 119.030 ;
        RECT 68.190 118.500 68.360 118.670 ;
        RECT 68.740 120.435 68.910 120.605 ;
        RECT 68.740 120.075 68.910 120.245 ;
        RECT 68.740 119.715 68.910 119.885 ;
        RECT 70.410 120.435 70.580 120.605 ;
        RECT 70.410 120.075 70.580 120.245 ;
        RECT 70.410 119.715 70.580 119.885 ;
        RECT 69.395 119.540 69.565 119.710 ;
        RECT 69.755 119.540 69.925 119.710 ;
        RECT 68.740 119.355 68.910 119.525 ;
        RECT 68.740 118.995 68.910 119.165 ;
        RECT 68.740 118.635 68.910 118.805 ;
        RECT 70.410 119.355 70.580 119.525 ;
        RECT 70.410 118.995 70.580 119.165 ;
        RECT 70.410 118.635 70.580 118.805 ;
        RECT 70.960 120.300 71.130 120.470 ;
        RECT 70.960 119.940 71.130 120.110 ;
        RECT 70.960 119.580 71.130 119.750 ;
        RECT 70.960 119.220 71.130 119.390 ;
        RECT 70.960 118.860 71.130 119.030 ;
        RECT 70.960 118.500 71.130 118.670 ;
        RECT 68.190 118.140 68.360 118.310 ;
        RECT 69.395 118.260 69.565 118.430 ;
        RECT 69.755 118.260 69.925 118.430 ;
        RECT 70.960 118.140 71.130 118.310 ;
        RECT 68.500 117.590 68.670 117.760 ;
        RECT 68.860 117.590 69.030 117.760 ;
        RECT 69.220 117.590 69.390 117.760 ;
        RECT 69.580 117.590 69.750 117.760 ;
        RECT 69.940 117.590 70.110 117.760 ;
        RECT 70.300 117.590 70.470 117.760 ;
        RECT 70.660 117.590 70.830 117.760 ;
        RECT 72.590 138.110 72.760 138.280 ;
        RECT 72.590 137.750 72.760 137.920 ;
        RECT 73.140 139.170 73.310 139.340 ;
        RECT 73.140 138.810 73.310 138.980 ;
        RECT 73.140 138.450 73.310 138.620 ;
        RECT 73.140 138.090 73.310 138.260 ;
        RECT 73.140 137.730 73.310 137.900 ;
        RECT 74.310 139.170 74.480 139.340 ;
        RECT 74.310 138.810 74.480 138.980 ;
        RECT 75.880 139.205 76.050 139.375 ;
        RECT 75.880 138.845 76.050 139.015 ;
        RECT 77.050 141.365 77.220 141.535 ;
        RECT 77.050 141.005 77.220 141.175 ;
        RECT 77.050 140.645 77.220 140.815 ;
        RECT 77.050 140.285 77.220 140.455 ;
        RECT 77.050 139.925 77.220 140.095 ;
        RECT 77.050 139.565 77.220 139.735 ;
        RECT 77.050 139.205 77.220 139.375 ;
        RECT 77.050 138.845 77.220 139.015 ;
        RECT 77.600 141.350 77.770 141.520 ;
        RECT 77.600 140.990 77.770 141.160 ;
        RECT 77.600 140.630 77.770 140.800 ;
        RECT 77.600 140.270 77.770 140.440 ;
        RECT 77.600 139.910 77.770 140.080 ;
        RECT 77.600 139.550 77.770 139.720 ;
        RECT 77.600 139.190 77.770 139.360 ;
        RECT 77.600 138.830 77.770 139.000 ;
        RECT 74.310 138.450 74.480 138.620 ;
        RECT 76.465 138.470 76.635 138.640 ;
        RECT 77.600 138.470 77.770 138.640 ;
        RECT 74.310 138.090 74.480 138.260 ;
        RECT 74.310 137.730 74.480 137.900 ;
        RECT 75.880 138.085 76.050 138.255 ;
        RECT 72.590 137.390 72.760 137.560 ;
        RECT 75.880 137.725 76.050 137.895 ;
        RECT 73.725 137.310 73.895 137.480 ;
        RECT 75.880 137.365 76.050 137.535 ;
        RECT 72.590 137.030 72.760 137.200 ;
        RECT 72.590 136.670 72.760 136.840 ;
        RECT 72.590 136.310 72.760 136.480 ;
        RECT 72.590 135.950 72.760 136.120 ;
        RECT 72.590 135.590 72.760 135.760 ;
        RECT 73.140 136.890 73.310 137.060 ;
        RECT 73.140 136.530 73.310 136.700 ;
        RECT 73.140 136.170 73.310 136.340 ;
        RECT 73.140 135.810 73.310 135.980 ;
        RECT 73.140 135.450 73.310 135.620 ;
        RECT 74.310 136.890 74.480 137.060 ;
        RECT 74.310 136.530 74.480 136.700 ;
        RECT 74.310 136.170 74.480 136.340 ;
        RECT 74.310 135.810 74.480 135.980 ;
        RECT 74.310 135.450 74.480 135.620 ;
        RECT 75.880 137.005 76.050 137.175 ;
        RECT 75.880 136.645 76.050 136.815 ;
        RECT 75.880 136.285 76.050 136.455 ;
        RECT 75.880 135.925 76.050 136.095 ;
        RECT 75.880 135.565 76.050 135.735 ;
        RECT 77.050 138.085 77.220 138.255 ;
        RECT 77.050 137.725 77.220 137.895 ;
        RECT 77.050 137.365 77.220 137.535 ;
        RECT 77.050 137.005 77.220 137.175 ;
        RECT 77.050 136.645 77.220 136.815 ;
        RECT 77.050 136.285 77.220 136.455 ;
        RECT 77.050 135.925 77.220 136.095 ;
        RECT 77.050 135.565 77.220 135.735 ;
        RECT 77.600 138.110 77.770 138.280 ;
        RECT 77.600 137.750 77.770 137.920 ;
        RECT 77.600 137.390 77.770 137.560 ;
        RECT 77.600 137.030 77.770 137.200 ;
        RECT 77.600 136.670 77.770 136.840 ;
        RECT 77.600 136.310 77.770 136.480 ;
        RECT 77.600 135.950 77.770 136.120 ;
        RECT 77.600 135.590 77.770 135.760 ;
        RECT 72.590 135.230 72.760 135.400 ;
        RECT 72.590 134.870 72.760 135.040 ;
        RECT 73.725 135.030 73.895 135.200 ;
        RECT 76.465 135.190 76.635 135.360 ;
        RECT 77.600 135.230 77.770 135.400 ;
        RECT 77.050 134.790 77.220 134.960 ;
        RECT 72.590 134.510 72.760 134.680 ;
        RECT 72.590 134.150 72.760 134.320 ;
        RECT 72.590 133.790 72.760 133.960 ;
        RECT 72.590 133.430 72.760 133.600 ;
        RECT 72.590 133.070 72.760 133.240 ;
        RECT 73.140 134.610 73.310 134.780 ;
        RECT 73.140 134.250 73.310 134.420 ;
        RECT 73.140 133.890 73.310 134.060 ;
        RECT 73.140 133.530 73.310 133.700 ;
        RECT 73.140 133.170 73.310 133.340 ;
        RECT 74.310 134.610 74.480 134.780 ;
        RECT 74.310 134.250 74.480 134.420 ;
        RECT 74.310 133.890 74.480 134.060 ;
        RECT 74.310 133.530 74.480 133.700 ;
        RECT 74.310 133.170 74.480 133.340 ;
        RECT 77.050 134.430 77.220 134.600 ;
        RECT 77.050 134.070 77.220 134.240 ;
        RECT 77.050 133.710 77.220 133.880 ;
        RECT 77.050 133.350 77.220 133.520 ;
        RECT 77.050 132.990 77.220 133.160 ;
        RECT 72.590 132.710 72.760 132.880 ;
        RECT 73.725 132.750 73.895 132.920 ;
        RECT 72.590 132.350 72.760 132.520 ;
        RECT 77.050 132.630 77.220 132.800 ;
        RECT 72.590 131.990 72.760 132.160 ;
        RECT 72.590 131.630 72.760 131.800 ;
        RECT 72.590 131.270 72.760 131.440 ;
        RECT 72.590 130.910 72.760 131.080 ;
        RECT 73.140 132.330 73.310 132.500 ;
        RECT 73.140 131.970 73.310 132.140 ;
        RECT 73.140 131.610 73.310 131.780 ;
        RECT 73.140 131.250 73.310 131.420 ;
        RECT 73.140 130.890 73.310 131.060 ;
        RECT 74.310 132.330 74.480 132.500 ;
        RECT 74.310 131.970 74.480 132.140 ;
        RECT 74.310 131.610 74.480 131.780 ;
        RECT 74.310 131.250 74.480 131.420 ;
        RECT 74.310 130.890 74.480 131.060 ;
        RECT 77.050 132.270 77.220 132.440 ;
        RECT 77.050 131.910 77.220 132.080 ;
        RECT 77.050 131.550 77.220 131.720 ;
        RECT 77.050 131.190 77.220 131.360 ;
        RECT 72.590 130.550 72.760 130.720 ;
        RECT 77.050 130.830 77.220 131.000 ;
        RECT 73.725 130.470 73.895 130.640 ;
        RECT 77.050 130.470 77.220 130.640 ;
        RECT 72.590 130.190 72.760 130.360 ;
        RECT 72.590 129.830 72.760 130.000 ;
        RECT 72.590 129.470 72.760 129.640 ;
        RECT 72.590 129.110 72.760 129.280 ;
        RECT 72.590 128.750 72.760 128.920 ;
        RECT 72.590 128.390 72.760 128.560 ;
        RECT 73.140 130.085 73.310 130.255 ;
        RECT 73.140 129.725 73.310 129.895 ;
        RECT 73.140 129.365 73.310 129.535 ;
        RECT 74.310 130.085 74.480 130.255 ;
        RECT 74.310 129.725 74.480 129.895 ;
        RECT 74.310 129.365 74.480 129.535 ;
        RECT 73.725 129.190 73.895 129.360 ;
        RECT 73.140 129.005 73.310 129.175 ;
        RECT 73.140 128.645 73.310 128.815 ;
        RECT 73.140 128.285 73.310 128.455 ;
        RECT 74.310 129.005 74.480 129.175 ;
        RECT 74.310 128.645 74.480 128.815 ;
        RECT 74.310 128.285 74.480 128.455 ;
        RECT 77.050 130.110 77.220 130.280 ;
        RECT 77.050 129.750 77.220 129.920 ;
        RECT 77.050 129.390 77.220 129.560 ;
        RECT 77.050 129.030 77.220 129.200 ;
        RECT 77.050 128.670 77.220 128.840 ;
        RECT 77.050 128.310 77.220 128.480 ;
        RECT 77.600 134.870 77.770 135.040 ;
        RECT 77.600 134.510 77.770 134.680 ;
        RECT 77.600 134.150 77.770 134.320 ;
        RECT 77.600 133.790 77.770 133.960 ;
        RECT 77.600 133.430 77.770 133.600 ;
        RECT 77.600 133.070 77.770 133.240 ;
        RECT 77.600 132.710 77.770 132.880 ;
        RECT 77.600 132.350 77.770 132.520 ;
        RECT 77.600 131.990 77.770 132.160 ;
        RECT 77.600 131.630 77.770 131.800 ;
        RECT 77.600 131.270 77.770 131.440 ;
        RECT 77.600 130.910 77.770 131.080 ;
        RECT 77.600 130.550 77.770 130.720 ;
        RECT 77.600 130.190 77.770 130.360 ;
        RECT 77.600 129.830 77.770 130.000 ;
        RECT 77.600 129.470 77.770 129.640 ;
        RECT 77.600 129.110 77.770 129.280 ;
        RECT 77.600 128.750 77.770 128.920 ;
        RECT 77.600 128.390 77.770 128.560 ;
        RECT 72.590 128.030 72.760 128.200 ;
        RECT 73.725 127.910 73.895 128.080 ;
        RECT 76.465 127.910 76.635 128.080 ;
        RECT 77.600 128.030 77.770 128.200 ;
        RECT 72.590 127.670 72.760 127.840 ;
        RECT 72.590 127.310 72.760 127.480 ;
        RECT 72.590 126.950 72.760 127.120 ;
        RECT 72.590 126.590 72.760 126.760 ;
        RECT 72.590 126.230 72.760 126.400 ;
        RECT 72.590 125.870 72.760 126.040 ;
        RECT 73.140 127.525 73.310 127.695 ;
        RECT 73.140 127.165 73.310 127.335 ;
        RECT 73.140 126.805 73.310 126.975 ;
        RECT 74.310 127.525 74.480 127.695 ;
        RECT 74.310 127.165 74.480 127.335 ;
        RECT 74.310 126.805 74.480 126.975 ;
        RECT 73.725 126.630 73.895 126.800 ;
        RECT 73.140 126.445 73.310 126.615 ;
        RECT 73.140 126.085 73.310 126.255 ;
        RECT 73.140 125.725 73.310 125.895 ;
        RECT 74.310 126.445 74.480 126.615 ;
        RECT 74.310 126.085 74.480 126.255 ;
        RECT 74.310 125.725 74.480 125.895 ;
        RECT 77.050 127.510 77.220 127.680 ;
        RECT 77.050 127.150 77.220 127.320 ;
        RECT 77.050 126.790 77.220 126.960 ;
        RECT 77.050 126.430 77.220 126.600 ;
        RECT 77.050 126.070 77.220 126.240 ;
        RECT 72.590 125.510 72.760 125.680 ;
        RECT 77.050 125.710 77.220 125.880 ;
        RECT 73.725 125.350 73.895 125.520 ;
        RECT 77.050 125.350 77.220 125.520 ;
        RECT 72.590 125.150 72.760 125.320 ;
        RECT 72.590 124.790 72.760 124.960 ;
        RECT 72.590 124.430 72.760 124.600 ;
        RECT 72.590 124.070 72.760 124.240 ;
        RECT 72.590 123.710 72.760 123.880 ;
        RECT 72.590 123.350 72.760 123.520 ;
        RECT 73.140 124.930 73.310 125.100 ;
        RECT 73.140 124.570 73.310 124.740 ;
        RECT 73.140 124.210 73.310 124.380 ;
        RECT 73.140 123.850 73.310 124.020 ;
        RECT 73.140 123.490 73.310 123.660 ;
        RECT 74.310 124.930 74.480 125.100 ;
        RECT 74.310 124.570 74.480 124.740 ;
        RECT 74.310 124.210 74.480 124.380 ;
        RECT 74.310 123.850 74.480 124.020 ;
        RECT 74.310 123.490 74.480 123.660 ;
        RECT 77.050 124.990 77.220 125.160 ;
        RECT 77.050 124.630 77.220 124.800 ;
        RECT 77.050 124.270 77.220 124.440 ;
        RECT 77.050 123.910 77.220 124.080 ;
        RECT 77.050 123.550 77.220 123.720 ;
        RECT 72.590 122.990 72.760 123.160 ;
        RECT 73.725 123.070 73.895 123.240 ;
        RECT 77.050 123.190 77.220 123.360 ;
        RECT 77.050 122.830 77.220 123.000 ;
        RECT 72.590 122.630 72.760 122.800 ;
        RECT 72.590 122.270 72.760 122.440 ;
        RECT 72.590 121.910 72.760 122.080 ;
        RECT 72.590 121.550 72.760 121.720 ;
        RECT 72.590 121.190 72.760 121.360 ;
        RECT 73.140 122.650 73.310 122.820 ;
        RECT 73.140 122.290 73.310 122.460 ;
        RECT 73.140 121.930 73.310 122.100 ;
        RECT 73.140 121.570 73.310 121.740 ;
        RECT 73.140 121.210 73.310 121.380 ;
        RECT 74.310 122.650 74.480 122.820 ;
        RECT 74.310 122.290 74.480 122.460 ;
        RECT 74.310 121.930 74.480 122.100 ;
        RECT 74.310 121.570 74.480 121.740 ;
        RECT 74.310 121.210 74.480 121.380 ;
        RECT 77.050 122.470 77.220 122.640 ;
        RECT 77.050 122.110 77.220 122.280 ;
        RECT 77.050 121.750 77.220 121.920 ;
        RECT 77.050 121.390 77.220 121.560 ;
        RECT 77.050 121.030 77.220 121.200 ;
        RECT 77.600 127.670 77.770 127.840 ;
        RECT 77.600 127.310 77.770 127.480 ;
        RECT 77.600 126.950 77.770 127.120 ;
        RECT 77.600 126.590 77.770 126.760 ;
        RECT 77.600 126.230 77.770 126.400 ;
        RECT 77.600 125.870 77.770 126.040 ;
        RECT 77.600 125.510 77.770 125.680 ;
        RECT 77.600 125.150 77.770 125.320 ;
        RECT 77.600 124.790 77.770 124.960 ;
        RECT 77.600 124.430 77.770 124.600 ;
        RECT 77.600 124.070 77.770 124.240 ;
        RECT 77.600 123.710 77.770 123.880 ;
        RECT 77.600 123.350 77.770 123.520 ;
        RECT 77.600 122.990 77.770 123.160 ;
        RECT 77.600 122.630 77.770 122.800 ;
        RECT 77.600 122.270 77.770 122.440 ;
        RECT 77.600 121.910 77.770 122.080 ;
        RECT 77.600 121.550 77.770 121.720 ;
        RECT 77.600 121.190 77.770 121.360 ;
        RECT 72.590 120.830 72.760 121.000 ;
        RECT 73.725 120.790 73.895 120.960 ;
        RECT 77.600 120.830 77.770 121.000 ;
        RECT 72.590 120.470 72.760 120.640 ;
        RECT 76.465 120.630 76.635 120.800 ;
        RECT 72.590 120.110 72.760 120.280 ;
        RECT 72.590 119.750 72.760 119.920 ;
        RECT 72.590 119.390 72.760 119.560 ;
        RECT 72.590 119.030 72.760 119.200 ;
        RECT 73.140 120.370 73.310 120.540 ;
        RECT 73.140 120.010 73.310 120.180 ;
        RECT 73.140 119.650 73.310 119.820 ;
        RECT 73.140 119.290 73.310 119.460 ;
        RECT 73.140 118.930 73.310 119.100 ;
        RECT 74.310 120.370 74.480 120.540 ;
        RECT 77.600 120.470 77.770 120.640 ;
        RECT 74.310 120.010 74.480 120.180 ;
        RECT 74.310 119.650 74.480 119.820 ;
        RECT 74.310 119.290 74.480 119.460 ;
        RECT 74.310 118.930 74.480 119.100 ;
        RECT 75.880 120.245 76.050 120.415 ;
        RECT 75.880 119.885 76.050 120.055 ;
        RECT 75.880 119.525 76.050 119.695 ;
        RECT 75.880 119.165 76.050 119.335 ;
        RECT 72.590 118.670 72.760 118.840 ;
        RECT 75.880 118.805 76.050 118.975 ;
        RECT 73.725 118.510 73.895 118.680 ;
        RECT 72.590 118.310 72.760 118.480 ;
        RECT 75.880 118.445 76.050 118.615 ;
        RECT 72.590 117.950 72.760 118.120 ;
        RECT 72.590 117.590 72.760 117.760 ;
        RECT 62.540 117.310 62.710 117.480 ;
        RECT 62.540 116.950 62.710 117.120 ;
        RECT 56.180 116.590 56.350 116.760 ;
        RECT 57.385 116.510 57.555 116.680 ;
        RECT 57.745 116.510 57.915 116.680 ;
        RECT 60.975 116.510 61.145 116.680 ;
        RECT 61.335 116.510 61.505 116.680 ;
        RECT 62.540 116.590 62.710 116.760 ;
        RECT 56.180 116.230 56.350 116.400 ;
        RECT 56.180 115.870 56.350 116.040 ;
        RECT 56.180 115.510 56.350 115.680 ;
        RECT 56.180 115.150 56.350 115.320 ;
        RECT 56.180 114.790 56.350 114.960 ;
        RECT 58.400 116.090 58.570 116.260 ;
        RECT 58.400 115.730 58.570 115.900 ;
        RECT 58.400 115.370 58.570 115.540 ;
        RECT 58.400 115.010 58.570 115.180 ;
        RECT 58.400 114.650 58.570 114.820 ;
        RECT 60.320 116.090 60.490 116.260 ;
        RECT 60.320 115.730 60.490 115.900 ;
        RECT 60.320 115.370 60.490 115.540 ;
        RECT 60.320 115.010 60.490 115.180 ;
        RECT 60.320 114.650 60.490 114.820 ;
        RECT 61.990 116.090 62.160 116.260 ;
        RECT 61.990 115.730 62.160 115.900 ;
        RECT 61.990 115.370 62.160 115.540 ;
        RECT 61.990 115.010 62.160 115.180 ;
        RECT 61.990 114.650 62.160 114.820 ;
        RECT 62.540 116.230 62.710 116.400 ;
        RECT 62.540 115.870 62.710 116.040 ;
        RECT 62.540 115.510 62.710 115.680 ;
        RECT 62.540 115.150 62.710 115.320 ;
        RECT 62.540 114.790 62.710 114.960 ;
        RECT 56.180 114.430 56.350 114.600 ;
        RECT 62.540 114.430 62.710 114.600 ;
        RECT 56.180 114.070 56.350 114.240 ;
        RECT 57.385 114.230 57.555 114.400 ;
        RECT 57.745 114.230 57.915 114.400 ;
        RECT 60.975 114.230 61.145 114.400 ;
        RECT 61.335 114.230 61.505 114.400 ;
        RECT 62.540 114.070 62.710 114.240 ;
        RECT 56.180 113.710 56.350 113.880 ;
        RECT 56.180 113.350 56.350 113.520 ;
        RECT 56.180 112.990 56.350 113.160 ;
        RECT 60.320 113.810 60.490 113.980 ;
        RECT 62.540 113.710 62.710 113.880 ;
        RECT 60.320 113.450 60.490 113.620 ;
        RECT 60.975 113.450 61.145 113.620 ;
        RECT 61.335 113.450 61.505 113.620 ;
        RECT 60.320 113.090 60.490 113.260 ;
        RECT 62.540 113.350 62.710 113.520 ;
        RECT 72.590 117.230 72.760 117.400 ;
        RECT 72.590 116.870 72.760 117.040 ;
        RECT 72.590 116.510 72.760 116.680 ;
        RECT 73.140 118.090 73.310 118.260 ;
        RECT 73.140 117.730 73.310 117.900 ;
        RECT 73.140 117.370 73.310 117.540 ;
        RECT 73.140 117.010 73.310 117.180 ;
        RECT 73.140 116.650 73.310 116.820 ;
        RECT 74.310 118.090 74.480 118.260 ;
        RECT 74.310 117.730 74.480 117.900 ;
        RECT 75.880 118.085 76.050 118.255 ;
        RECT 75.880 117.725 76.050 117.895 ;
        RECT 77.050 120.245 77.220 120.415 ;
        RECT 77.050 119.885 77.220 120.055 ;
        RECT 77.050 119.525 77.220 119.695 ;
        RECT 77.050 119.165 77.220 119.335 ;
        RECT 77.050 118.805 77.220 118.975 ;
        RECT 77.050 118.445 77.220 118.615 ;
        RECT 77.050 118.085 77.220 118.255 ;
        RECT 77.050 117.725 77.220 117.895 ;
        RECT 77.600 120.110 77.770 120.280 ;
        RECT 77.600 119.750 77.770 119.920 ;
        RECT 77.600 119.390 77.770 119.560 ;
        RECT 77.600 119.030 77.770 119.200 ;
        RECT 77.600 118.670 77.770 118.840 ;
        RECT 77.600 118.310 77.770 118.480 ;
        RECT 77.600 117.950 77.770 118.120 ;
        RECT 74.310 117.370 74.480 117.540 ;
        RECT 77.600 117.590 77.770 117.760 ;
        RECT 76.465 117.350 76.635 117.520 ;
        RECT 74.310 117.010 74.480 117.180 ;
        RECT 77.600 117.230 77.770 117.400 ;
        RECT 74.310 116.650 74.480 116.820 ;
        RECT 75.880 116.965 76.050 117.135 ;
        RECT 75.880 116.605 76.050 116.775 ;
        RECT 72.590 116.150 72.760 116.320 ;
        RECT 73.725 116.230 73.895 116.400 ;
        RECT 75.880 116.245 76.050 116.415 ;
        RECT 72.590 115.790 72.760 115.960 ;
        RECT 72.590 115.430 72.760 115.600 ;
        RECT 72.590 115.070 72.760 115.240 ;
        RECT 74.310 115.845 74.480 116.015 ;
        RECT 74.310 115.485 74.480 115.655 ;
        RECT 74.310 115.125 74.480 115.295 ;
        RECT 73.725 114.950 73.895 115.120 ;
        RECT 72.590 114.710 72.760 114.880 ;
        RECT 72.590 114.350 72.760 114.520 ;
        RECT 72.590 113.990 72.760 114.160 ;
        RECT 74.310 114.765 74.480 114.935 ;
        RECT 74.310 114.405 74.480 114.575 ;
        RECT 75.880 115.885 76.050 116.055 ;
        RECT 75.880 115.525 76.050 115.695 ;
        RECT 75.880 115.165 76.050 115.335 ;
        RECT 75.880 114.805 76.050 114.975 ;
        RECT 75.880 114.445 76.050 114.615 ;
        RECT 77.050 116.965 77.220 117.135 ;
        RECT 77.050 116.605 77.220 116.775 ;
        RECT 77.050 116.245 77.220 116.415 ;
        RECT 77.050 115.885 77.220 116.055 ;
        RECT 77.050 115.525 77.220 115.695 ;
        RECT 77.050 115.165 77.220 115.335 ;
        RECT 77.050 114.805 77.220 114.975 ;
        RECT 77.050 114.445 77.220 114.615 ;
        RECT 77.600 116.870 77.770 117.040 ;
        RECT 77.600 116.510 77.770 116.680 ;
        RECT 77.600 116.150 77.770 116.320 ;
        RECT 77.600 115.790 77.770 115.960 ;
        RECT 77.600 115.430 77.770 115.600 ;
        RECT 77.600 115.070 77.770 115.240 ;
        RECT 77.600 114.710 77.770 114.880 ;
        RECT 77.600 114.350 77.770 114.520 ;
        RECT 74.310 114.045 74.480 114.215 ;
        RECT 76.465 114.070 76.635 114.240 ;
        RECT 77.600 113.990 77.770 114.160 ;
        RECT 72.590 113.630 72.760 113.800 ;
        RECT 73.725 113.670 73.895 113.840 ;
        RECT 62.540 112.990 62.710 113.160 ;
        RECT 56.180 112.630 56.350 112.800 ;
        RECT 60.975 112.670 61.145 112.840 ;
        RECT 61.335 112.670 61.505 112.840 ;
        RECT 62.540 112.630 62.710 112.800 ;
        RECT 56.480 112.000 56.650 112.170 ;
        RECT 56.840 112.000 57.010 112.170 ;
        RECT 57.200 112.000 57.370 112.170 ;
        RECT 57.560 112.000 57.730 112.170 ;
        RECT 57.920 112.000 58.090 112.170 ;
        RECT 58.280 112.000 58.450 112.170 ;
        RECT 58.640 112.000 58.810 112.170 ;
        RECT 59.000 112.000 59.170 112.170 ;
        RECT 59.360 112.000 59.530 112.170 ;
        RECT 59.720 112.000 59.890 112.170 ;
        RECT 60.080 112.000 60.250 112.170 ;
        RECT 60.440 112.000 60.610 112.170 ;
        RECT 60.800 112.000 60.970 112.170 ;
        RECT 61.160 112.000 61.330 112.170 ;
        RECT 61.520 112.000 61.690 112.170 ;
        RECT 61.880 112.000 62.050 112.170 ;
        RECT 62.240 112.000 62.410 112.170 ;
        RECT 63.985 113.340 64.155 113.510 ;
        RECT 64.345 113.340 64.515 113.510 ;
        RECT 64.705 113.340 64.875 113.510 ;
        RECT 65.065 113.340 65.235 113.510 ;
        RECT 65.425 113.340 65.595 113.510 ;
        RECT 65.785 113.340 65.955 113.510 ;
        RECT 66.145 113.340 66.315 113.510 ;
        RECT 66.505 113.340 66.675 113.510 ;
        RECT 67.975 113.340 68.145 113.510 ;
        RECT 68.335 113.340 68.505 113.510 ;
        RECT 68.695 113.340 68.865 113.510 ;
        RECT 69.055 113.340 69.225 113.510 ;
        RECT 69.415 113.340 69.585 113.510 ;
        RECT 69.775 113.340 69.945 113.510 ;
        RECT 63.685 112.990 63.855 113.160 ;
        RECT 70.075 112.990 70.245 113.160 ;
        RECT 77.600 113.630 77.770 113.800 ;
        RECT 72.980 113.040 73.150 113.210 ;
        RECT 73.340 113.040 73.510 113.210 ;
        RECT 73.700 113.040 73.870 113.210 ;
        RECT 74.060 113.040 74.230 113.210 ;
        RECT 74.420 113.040 74.590 113.210 ;
        RECT 74.780 113.040 74.950 113.210 ;
        RECT 75.140 113.040 75.310 113.210 ;
        RECT 75.500 113.040 75.670 113.210 ;
        RECT 75.860 113.040 76.030 113.210 ;
        RECT 76.220 113.040 76.390 113.210 ;
        RECT 76.580 113.040 76.750 113.210 ;
        RECT 76.940 113.040 77.110 113.210 ;
        RECT 77.300 113.040 77.470 113.210 ;
        RECT 81.320 142.780 81.490 142.950 ;
        RECT 81.680 142.780 81.850 142.950 ;
        RECT 82.040 142.780 82.210 142.950 ;
        RECT 82.400 142.780 82.570 142.950 ;
        RECT 82.760 142.780 82.930 142.950 ;
        RECT 83.120 142.780 83.290 142.950 ;
        RECT 83.480 142.780 83.650 142.950 ;
        RECT 83.840 142.780 84.010 142.950 ;
        RECT 84.200 142.780 84.370 142.950 ;
        RECT 84.560 142.780 84.730 142.950 ;
        RECT 84.920 142.780 85.090 142.950 ;
        RECT 85.280 142.780 85.450 142.950 ;
        RECT 85.640 142.780 85.810 142.950 ;
        RECT 81.020 142.430 81.190 142.600 ;
        RECT 86.030 142.430 86.200 142.600 ;
        RECT 91.915 142.870 92.085 143.040 ;
        RECT 94.185 142.870 94.355 143.040 ;
        RECT 92.215 142.480 92.385 142.650 ;
        RECT 92.575 142.480 92.745 142.650 ;
        RECT 92.935 142.480 93.105 142.650 ;
        RECT 93.295 142.480 93.465 142.650 ;
        RECT 93.655 142.480 93.825 142.650 ;
        RECT 96.380 151.500 96.550 151.670 ;
        RECT 96.740 151.500 96.910 151.670 ;
        RECT 97.100 151.500 97.270 151.670 ;
        RECT 97.460 151.500 97.630 151.670 ;
        RECT 97.820 151.500 97.990 151.670 ;
        RECT 98.180 151.500 98.350 151.670 ;
        RECT 98.540 151.500 98.710 151.670 ;
        RECT 98.900 151.500 99.070 151.670 ;
        RECT 99.260 151.500 99.430 151.670 ;
        RECT 99.620 151.500 99.790 151.670 ;
        RECT 99.980 151.500 100.150 151.670 ;
        RECT 100.340 151.500 100.510 151.670 ;
        RECT 100.700 151.500 100.870 151.670 ;
        RECT 101.060 151.500 101.230 151.670 ;
        RECT 101.420 151.500 101.590 151.670 ;
        RECT 101.780 151.500 101.950 151.670 ;
        RECT 102.140 151.500 102.310 151.670 ;
        RECT 96.080 151.150 96.250 151.320 ;
        RECT 102.440 151.150 102.610 151.320 ;
        RECT 96.080 150.790 96.250 150.960 ;
        RECT 97.285 150.830 97.455 151.000 ;
        RECT 97.645 150.830 97.815 151.000 ;
        RECT 96.080 150.430 96.250 150.600 ;
        RECT 102.440 150.790 102.610 150.960 ;
        RECT 96.080 150.070 96.250 150.240 ;
        RECT 98.300 150.410 98.470 150.580 ;
        RECT 97.285 150.050 97.455 150.220 ;
        RECT 97.645 150.050 97.815 150.220 ;
        RECT 98.300 150.050 98.470 150.220 ;
        RECT 96.080 149.710 96.250 149.880 ;
        RECT 98.300 149.690 98.470 149.860 ;
        RECT 102.440 150.430 102.610 150.600 ;
        RECT 102.440 150.070 102.610 150.240 ;
        RECT 102.440 149.710 102.610 149.880 ;
        RECT 96.080 149.350 96.250 149.520 ;
        RECT 97.285 149.270 97.455 149.440 ;
        RECT 97.645 149.270 97.815 149.440 ;
        RECT 102.440 149.350 102.610 149.520 ;
        RECT 96.080 148.990 96.250 149.160 ;
        RECT 96.080 148.630 96.250 148.800 ;
        RECT 96.080 148.270 96.250 148.440 ;
        RECT 96.080 147.910 96.250 148.080 ;
        RECT 96.080 147.550 96.250 147.720 ;
        RECT 96.630 148.850 96.800 149.020 ;
        RECT 96.630 148.490 96.800 148.660 ;
        RECT 96.630 148.130 96.800 148.300 ;
        RECT 96.630 147.770 96.800 147.940 ;
        RECT 96.630 147.410 96.800 147.580 ;
        RECT 102.440 148.990 102.610 149.160 ;
        RECT 102.440 148.630 102.610 148.800 ;
        RECT 102.440 148.270 102.610 148.440 ;
        RECT 102.440 147.910 102.610 148.080 ;
        RECT 102.440 147.550 102.610 147.720 ;
        RECT 96.080 147.190 96.250 147.360 ;
        RECT 102.440 147.190 102.610 147.360 ;
        RECT 96.080 146.830 96.250 147.000 ;
        RECT 97.285 146.990 97.455 147.160 ;
        RECT 97.645 146.990 97.815 147.160 ;
        RECT 102.440 146.830 102.610 147.000 ;
        RECT 96.080 146.470 96.250 146.640 ;
        RECT 96.080 146.110 96.250 146.280 ;
        RECT 96.080 145.750 96.250 145.920 ;
        RECT 96.080 145.390 96.250 145.560 ;
        RECT 96.080 145.030 96.250 145.200 ;
        RECT 96.630 146.570 96.800 146.740 ;
        RECT 96.630 146.210 96.800 146.380 ;
        RECT 96.630 145.850 96.800 146.020 ;
        RECT 96.630 145.490 96.800 145.660 ;
        RECT 96.630 145.130 96.800 145.300 ;
        RECT 102.440 146.470 102.610 146.640 ;
        RECT 102.440 146.110 102.610 146.280 ;
        RECT 102.440 145.750 102.610 145.920 ;
        RECT 102.440 145.390 102.610 145.560 ;
        RECT 102.440 145.030 102.610 145.200 ;
        RECT 96.080 144.670 96.250 144.840 ;
        RECT 97.285 144.710 97.455 144.880 ;
        RECT 97.645 144.710 97.815 144.880 ;
        RECT 96.080 144.310 96.250 144.480 ;
        RECT 102.440 144.670 102.610 144.840 ;
        RECT 96.080 143.950 96.250 144.120 ;
        RECT 98.300 144.290 98.470 144.460 ;
        RECT 97.285 143.930 97.455 144.100 ;
        RECT 97.645 143.930 97.815 144.100 ;
        RECT 98.300 143.930 98.470 144.100 ;
        RECT 96.080 143.590 96.250 143.760 ;
        RECT 98.300 143.570 98.470 143.740 ;
        RECT 102.440 144.310 102.610 144.480 ;
        RECT 102.440 143.950 102.610 144.120 ;
        RECT 102.440 143.590 102.610 143.760 ;
        RECT 96.080 143.230 96.250 143.400 ;
        RECT 97.285 143.150 97.455 143.320 ;
        RECT 97.645 143.150 97.815 143.320 ;
        RECT 102.440 143.230 102.610 143.400 ;
        RECT 96.080 142.870 96.250 143.040 ;
        RECT 96.080 142.510 96.250 142.680 ;
        RECT 98.300 142.730 98.470 142.900 ;
        RECT 81.020 142.070 81.190 142.240 ;
        RECT 84.895 142.150 85.065 142.320 ;
        RECT 86.030 142.070 86.200 142.240 ;
        RECT 81.020 141.710 81.190 141.880 ;
        RECT 82.155 141.750 82.325 141.920 ;
        RECT 84.310 141.765 84.480 141.935 ;
        RECT 81.020 141.350 81.190 141.520 ;
        RECT 81.020 140.990 81.190 141.160 ;
        RECT 81.020 140.630 81.190 140.800 ;
        RECT 81.020 140.270 81.190 140.440 ;
        RECT 81.020 139.910 81.190 140.080 ;
        RECT 81.020 139.550 81.190 139.720 ;
        RECT 81.020 139.190 81.190 139.360 ;
        RECT 81.020 138.830 81.190 139.000 ;
        RECT 81.570 141.365 81.740 141.535 ;
        RECT 81.570 141.005 81.740 141.175 ;
        RECT 81.570 140.645 81.740 140.815 ;
        RECT 81.570 140.285 81.740 140.455 ;
        RECT 81.570 139.925 81.740 140.095 ;
        RECT 81.570 139.565 81.740 139.735 ;
        RECT 81.570 139.205 81.740 139.375 ;
        RECT 81.570 138.845 81.740 139.015 ;
        RECT 82.740 141.365 82.910 141.535 ;
        RECT 82.740 141.005 82.910 141.175 ;
        RECT 82.740 140.645 82.910 140.815 ;
        RECT 82.740 140.285 82.910 140.455 ;
        RECT 82.740 139.925 82.910 140.095 ;
        RECT 84.310 141.405 84.480 141.575 ;
        RECT 84.310 141.045 84.480 141.215 ;
        RECT 86.030 141.710 86.200 141.880 ;
        RECT 86.030 141.350 86.200 141.520 ;
        RECT 84.895 140.870 85.065 141.040 ;
        RECT 86.030 140.990 86.200 141.160 ;
        RECT 84.310 140.685 84.480 140.855 ;
        RECT 84.310 140.325 84.480 140.495 ;
        RECT 84.310 139.965 84.480 140.135 ;
        RECT 86.030 140.630 86.200 140.800 ;
        RECT 86.030 140.270 86.200 140.440 ;
        RECT 86.030 139.910 86.200 140.080 ;
        RECT 82.740 139.565 82.910 139.735 ;
        RECT 84.895 139.590 85.065 139.760 ;
        RECT 82.740 139.205 82.910 139.375 ;
        RECT 86.030 139.550 86.200 139.720 ;
        RECT 82.740 138.845 82.910 139.015 ;
        RECT 84.310 139.170 84.480 139.340 ;
        RECT 84.310 138.810 84.480 138.980 ;
        RECT 81.020 138.470 81.190 138.640 ;
        RECT 82.155 138.470 82.325 138.640 ;
        RECT 81.020 138.110 81.190 138.280 ;
        RECT 84.310 138.450 84.480 138.620 ;
        RECT 81.020 137.750 81.190 137.920 ;
        RECT 81.020 137.390 81.190 137.560 ;
        RECT 81.020 137.030 81.190 137.200 ;
        RECT 81.020 136.670 81.190 136.840 ;
        RECT 81.020 136.310 81.190 136.480 ;
        RECT 81.020 135.950 81.190 136.120 ;
        RECT 81.020 135.590 81.190 135.760 ;
        RECT 81.570 138.085 81.740 138.255 ;
        RECT 81.570 137.725 81.740 137.895 ;
        RECT 81.570 137.365 81.740 137.535 ;
        RECT 81.570 137.005 81.740 137.175 ;
        RECT 81.570 136.645 81.740 136.815 ;
        RECT 81.570 136.285 81.740 136.455 ;
        RECT 81.570 135.925 81.740 136.095 ;
        RECT 81.570 135.565 81.740 135.735 ;
        RECT 82.740 138.085 82.910 138.255 ;
        RECT 82.740 137.725 82.910 137.895 ;
        RECT 84.310 138.090 84.480 138.260 ;
        RECT 84.310 137.730 84.480 137.900 ;
        RECT 85.480 139.170 85.650 139.340 ;
        RECT 85.480 138.810 85.650 138.980 ;
        RECT 85.480 138.450 85.650 138.620 ;
        RECT 85.480 138.090 85.650 138.260 ;
        RECT 85.480 137.730 85.650 137.900 ;
        RECT 86.030 139.190 86.200 139.360 ;
        RECT 86.030 138.830 86.200 139.000 ;
        RECT 86.030 138.470 86.200 138.640 ;
        RECT 97.285 142.370 97.455 142.540 ;
        RECT 97.645 142.370 97.815 142.540 ;
        RECT 98.300 142.370 98.470 142.540 ;
        RECT 96.080 142.150 96.250 142.320 ;
        RECT 98.300 142.010 98.470 142.180 ;
        RECT 102.440 142.870 102.610 143.040 ;
        RECT 102.440 142.510 102.610 142.680 ;
        RECT 102.440 142.150 102.610 142.320 ;
        RECT 96.080 141.790 96.250 141.960 ;
        RECT 102.440 141.790 102.610 141.960 ;
        RECT 96.080 141.430 96.250 141.600 ;
        RECT 97.285 141.590 97.455 141.760 ;
        RECT 97.645 141.590 97.815 141.760 ;
        RECT 100.875 141.590 101.045 141.760 ;
        RECT 101.235 141.590 101.405 141.760 ;
        RECT 102.440 141.430 102.610 141.600 ;
        RECT 96.080 141.070 96.250 141.240 ;
        RECT 96.080 140.710 96.250 140.880 ;
        RECT 96.080 140.350 96.250 140.520 ;
        RECT 96.080 139.990 96.250 140.160 ;
        RECT 96.080 139.630 96.250 139.800 ;
        RECT 96.630 141.170 96.800 141.340 ;
        RECT 96.630 140.810 96.800 140.980 ;
        RECT 96.630 140.450 96.800 140.620 ;
        RECT 96.630 140.090 96.800 140.260 ;
        RECT 96.630 139.730 96.800 139.900 ;
        RECT 98.300 141.170 98.470 141.340 ;
        RECT 98.300 140.810 98.470 140.980 ;
        RECT 98.300 140.450 98.470 140.620 ;
        RECT 98.300 140.090 98.470 140.260 ;
        RECT 98.300 139.730 98.470 139.900 ;
        RECT 100.220 141.170 100.390 141.340 ;
        RECT 100.220 140.810 100.390 140.980 ;
        RECT 100.220 140.450 100.390 140.620 ;
        RECT 100.220 140.090 100.390 140.260 ;
        RECT 100.220 139.730 100.390 139.900 ;
        RECT 102.440 141.070 102.610 141.240 ;
        RECT 102.440 140.710 102.610 140.880 ;
        RECT 102.440 140.350 102.610 140.520 ;
        RECT 102.440 139.990 102.610 140.160 ;
        RECT 102.440 139.630 102.610 139.800 ;
        RECT 96.080 139.270 96.250 139.440 ;
        RECT 97.285 139.310 97.455 139.480 ;
        RECT 97.645 139.310 97.815 139.480 ;
        RECT 100.875 139.310 101.045 139.480 ;
        RECT 101.235 139.310 101.405 139.480 ;
        RECT 96.080 138.910 96.250 139.080 ;
        RECT 102.440 139.270 102.610 139.440 ;
        RECT 96.080 138.550 96.250 138.720 ;
        RECT 86.030 138.110 86.200 138.280 ;
        RECT 86.030 137.750 86.200 137.920 ;
        RECT 82.740 137.365 82.910 137.535 ;
        RECT 84.895 137.310 85.065 137.480 ;
        RECT 86.030 137.390 86.200 137.560 ;
        RECT 82.740 137.005 82.910 137.175 ;
        RECT 82.740 136.645 82.910 136.815 ;
        RECT 82.740 136.285 82.910 136.455 ;
        RECT 82.740 135.925 82.910 136.095 ;
        RECT 82.740 135.565 82.910 135.735 ;
        RECT 84.310 136.890 84.480 137.060 ;
        RECT 84.310 136.530 84.480 136.700 ;
        RECT 84.310 136.170 84.480 136.340 ;
        RECT 84.310 135.810 84.480 135.980 ;
        RECT 84.310 135.450 84.480 135.620 ;
        RECT 85.480 136.890 85.650 137.060 ;
        RECT 85.480 136.530 85.650 136.700 ;
        RECT 85.480 136.170 85.650 136.340 ;
        RECT 85.480 135.810 85.650 135.980 ;
        RECT 85.480 135.450 85.650 135.620 ;
        RECT 86.030 137.030 86.200 137.200 ;
        RECT 86.030 136.670 86.200 136.840 ;
        RECT 86.030 136.310 86.200 136.480 ;
        RECT 86.030 135.950 86.200 136.120 ;
        RECT 86.030 135.590 86.200 135.760 ;
        RECT 81.020 135.230 81.190 135.400 ;
        RECT 82.155 135.190 82.325 135.360 ;
        RECT 86.030 135.230 86.200 135.400 ;
        RECT 81.020 134.870 81.190 135.040 ;
        RECT 84.895 135.030 85.065 135.200 ;
        RECT 81.020 134.510 81.190 134.680 ;
        RECT 81.020 134.150 81.190 134.320 ;
        RECT 81.020 133.790 81.190 133.960 ;
        RECT 81.020 133.430 81.190 133.600 ;
        RECT 81.020 133.070 81.190 133.240 ;
        RECT 81.020 132.710 81.190 132.880 ;
        RECT 81.020 132.350 81.190 132.520 ;
        RECT 81.020 131.990 81.190 132.160 ;
        RECT 81.020 131.630 81.190 131.800 ;
        RECT 81.020 131.270 81.190 131.440 ;
        RECT 81.020 130.910 81.190 131.080 ;
        RECT 81.020 130.550 81.190 130.720 ;
        RECT 81.020 130.190 81.190 130.360 ;
        RECT 81.020 129.830 81.190 130.000 ;
        RECT 81.020 129.470 81.190 129.640 ;
        RECT 81.020 129.110 81.190 129.280 ;
        RECT 81.020 128.750 81.190 128.920 ;
        RECT 81.020 128.390 81.190 128.560 ;
        RECT 81.570 134.790 81.740 134.960 ;
        RECT 86.030 134.870 86.200 135.040 ;
        RECT 81.570 134.430 81.740 134.600 ;
        RECT 81.570 134.070 81.740 134.240 ;
        RECT 81.570 133.710 81.740 133.880 ;
        RECT 81.570 133.350 81.740 133.520 ;
        RECT 84.310 134.610 84.480 134.780 ;
        RECT 84.310 134.250 84.480 134.420 ;
        RECT 84.310 133.890 84.480 134.060 ;
        RECT 84.310 133.530 84.480 133.700 ;
        RECT 84.310 133.170 84.480 133.340 ;
        RECT 85.480 134.610 85.650 134.780 ;
        RECT 85.480 134.250 85.650 134.420 ;
        RECT 85.480 133.890 85.650 134.060 ;
        RECT 85.480 133.530 85.650 133.700 ;
        RECT 85.480 133.170 85.650 133.340 ;
        RECT 86.030 134.510 86.200 134.680 ;
        RECT 86.030 134.150 86.200 134.320 ;
        RECT 86.030 133.790 86.200 133.960 ;
        RECT 86.030 133.430 86.200 133.600 ;
        RECT 81.570 132.990 81.740 133.160 ;
        RECT 86.030 133.070 86.200 133.240 ;
        RECT 81.570 132.630 81.740 132.800 ;
        RECT 84.895 132.750 85.065 132.920 ;
        RECT 86.030 132.710 86.200 132.880 ;
        RECT 81.570 132.270 81.740 132.440 ;
        RECT 81.570 131.910 81.740 132.080 ;
        RECT 81.570 131.550 81.740 131.720 ;
        RECT 81.570 131.190 81.740 131.360 ;
        RECT 81.570 130.830 81.740 131.000 ;
        RECT 84.310 132.330 84.480 132.500 ;
        RECT 84.310 131.970 84.480 132.140 ;
        RECT 84.310 131.610 84.480 131.780 ;
        RECT 84.310 131.250 84.480 131.420 ;
        RECT 84.310 130.890 84.480 131.060 ;
        RECT 85.480 132.330 85.650 132.500 ;
        RECT 85.480 131.970 85.650 132.140 ;
        RECT 85.480 131.610 85.650 131.780 ;
        RECT 85.480 131.250 85.650 131.420 ;
        RECT 85.480 130.890 85.650 131.060 ;
        RECT 86.030 132.350 86.200 132.520 ;
        RECT 86.030 131.990 86.200 132.160 ;
        RECT 86.030 131.630 86.200 131.800 ;
        RECT 86.030 131.270 86.200 131.440 ;
        RECT 86.030 130.910 86.200 131.080 ;
        RECT 81.570 130.470 81.740 130.640 ;
        RECT 84.895 130.470 85.065 130.640 ;
        RECT 86.030 130.550 86.200 130.720 ;
        RECT 81.570 130.110 81.740 130.280 ;
        RECT 81.570 129.750 81.740 129.920 ;
        RECT 81.570 129.390 81.740 129.560 ;
        RECT 81.570 129.030 81.740 129.200 ;
        RECT 81.570 128.670 81.740 128.840 ;
        RECT 81.570 128.310 81.740 128.480 ;
        RECT 84.310 130.085 84.480 130.255 ;
        RECT 84.310 129.725 84.480 129.895 ;
        RECT 84.310 129.365 84.480 129.535 ;
        RECT 85.480 130.085 85.650 130.255 ;
        RECT 85.480 129.725 85.650 129.895 ;
        RECT 85.480 129.365 85.650 129.535 ;
        RECT 84.895 129.190 85.065 129.360 ;
        RECT 84.310 129.005 84.480 129.175 ;
        RECT 84.310 128.645 84.480 128.815 ;
        RECT 84.310 128.285 84.480 128.455 ;
        RECT 85.480 129.005 85.650 129.175 ;
        RECT 85.480 128.645 85.650 128.815 ;
        RECT 85.480 128.285 85.650 128.455 ;
        RECT 86.030 130.190 86.200 130.360 ;
        RECT 86.030 129.830 86.200 130.000 ;
        RECT 86.030 129.470 86.200 129.640 ;
        RECT 86.030 129.110 86.200 129.280 ;
        RECT 86.030 128.750 86.200 128.920 ;
        RECT 86.030 128.390 86.200 128.560 ;
        RECT 81.020 128.030 81.190 128.200 ;
        RECT 82.155 127.910 82.325 128.080 ;
        RECT 84.895 127.910 85.065 128.080 ;
        RECT 86.030 128.030 86.200 128.200 ;
        RECT 81.020 127.670 81.190 127.840 ;
        RECT 81.020 127.310 81.190 127.480 ;
        RECT 81.020 126.950 81.190 127.120 ;
        RECT 81.020 126.590 81.190 126.760 ;
        RECT 81.020 126.230 81.190 126.400 ;
        RECT 81.020 125.870 81.190 126.040 ;
        RECT 81.020 125.510 81.190 125.680 ;
        RECT 81.020 125.150 81.190 125.320 ;
        RECT 81.020 124.790 81.190 124.960 ;
        RECT 81.020 124.430 81.190 124.600 ;
        RECT 81.020 124.070 81.190 124.240 ;
        RECT 81.020 123.710 81.190 123.880 ;
        RECT 81.020 123.350 81.190 123.520 ;
        RECT 81.020 122.990 81.190 123.160 ;
        RECT 81.020 122.630 81.190 122.800 ;
        RECT 81.020 122.270 81.190 122.440 ;
        RECT 81.020 121.910 81.190 122.080 ;
        RECT 81.020 121.550 81.190 121.720 ;
        RECT 81.020 121.190 81.190 121.360 ;
        RECT 81.570 127.510 81.740 127.680 ;
        RECT 81.570 127.150 81.740 127.320 ;
        RECT 81.570 126.790 81.740 126.960 ;
        RECT 81.570 126.430 81.740 126.600 ;
        RECT 81.570 126.070 81.740 126.240 ;
        RECT 81.570 125.710 81.740 125.880 ;
        RECT 84.310 127.525 84.480 127.695 ;
        RECT 84.310 127.165 84.480 127.335 ;
        RECT 84.310 126.805 84.480 126.975 ;
        RECT 85.480 127.525 85.650 127.695 ;
        RECT 85.480 127.165 85.650 127.335 ;
        RECT 85.480 126.805 85.650 126.975 ;
        RECT 84.895 126.630 85.065 126.800 ;
        RECT 84.310 126.445 84.480 126.615 ;
        RECT 84.310 126.085 84.480 126.255 ;
        RECT 84.310 125.725 84.480 125.895 ;
        RECT 85.480 126.445 85.650 126.615 ;
        RECT 85.480 126.085 85.650 126.255 ;
        RECT 85.480 125.725 85.650 125.895 ;
        RECT 86.030 127.670 86.200 127.840 ;
        RECT 86.030 127.310 86.200 127.480 ;
        RECT 86.030 126.950 86.200 127.120 ;
        RECT 86.030 126.590 86.200 126.760 ;
        RECT 86.030 126.230 86.200 126.400 ;
        RECT 86.030 125.870 86.200 126.040 ;
        RECT 81.570 125.350 81.740 125.520 ;
        RECT 84.895 125.350 85.065 125.520 ;
        RECT 86.030 125.510 86.200 125.680 ;
        RECT 81.570 124.990 81.740 125.160 ;
        RECT 86.030 125.150 86.200 125.320 ;
        RECT 81.570 124.630 81.740 124.800 ;
        RECT 81.570 124.270 81.740 124.440 ;
        RECT 81.570 123.910 81.740 124.080 ;
        RECT 81.570 123.550 81.740 123.720 ;
        RECT 84.310 124.930 84.480 125.100 ;
        RECT 84.310 124.570 84.480 124.740 ;
        RECT 84.310 124.210 84.480 124.380 ;
        RECT 84.310 123.850 84.480 124.020 ;
        RECT 84.310 123.490 84.480 123.660 ;
        RECT 85.480 124.930 85.650 125.100 ;
        RECT 85.480 124.570 85.650 124.740 ;
        RECT 85.480 124.210 85.650 124.380 ;
        RECT 85.480 123.850 85.650 124.020 ;
        RECT 85.480 123.490 85.650 123.660 ;
        RECT 86.030 124.790 86.200 124.960 ;
        RECT 86.030 124.430 86.200 124.600 ;
        RECT 86.030 124.070 86.200 124.240 ;
        RECT 86.030 123.710 86.200 123.880 ;
        RECT 81.570 123.190 81.740 123.360 ;
        RECT 86.030 123.350 86.200 123.520 ;
        RECT 84.895 123.070 85.065 123.240 ;
        RECT 81.570 122.830 81.740 123.000 ;
        RECT 86.030 122.990 86.200 123.160 ;
        RECT 81.570 122.470 81.740 122.640 ;
        RECT 81.570 122.110 81.740 122.280 ;
        RECT 81.570 121.750 81.740 121.920 ;
        RECT 81.570 121.390 81.740 121.560 ;
        RECT 84.310 122.650 84.480 122.820 ;
        RECT 84.310 122.290 84.480 122.460 ;
        RECT 84.310 121.930 84.480 122.100 ;
        RECT 84.310 121.570 84.480 121.740 ;
        RECT 84.310 121.210 84.480 121.380 ;
        RECT 85.480 122.650 85.650 122.820 ;
        RECT 85.480 122.290 85.650 122.460 ;
        RECT 85.480 121.930 85.650 122.100 ;
        RECT 85.480 121.570 85.650 121.740 ;
        RECT 85.480 121.210 85.650 121.380 ;
        RECT 86.030 122.630 86.200 122.800 ;
        RECT 86.030 122.270 86.200 122.440 ;
        RECT 86.030 121.910 86.200 122.080 ;
        RECT 86.030 121.550 86.200 121.720 ;
        RECT 81.570 121.030 81.740 121.200 ;
        RECT 86.030 121.190 86.200 121.360 ;
        RECT 81.020 120.830 81.190 121.000 ;
        RECT 81.020 120.470 81.190 120.640 ;
        RECT 82.155 120.630 82.325 120.800 ;
        RECT 84.895 120.790 85.065 120.960 ;
        RECT 86.030 120.830 86.200 121.000 ;
        RECT 81.020 120.110 81.190 120.280 ;
        RECT 81.020 119.750 81.190 119.920 ;
        RECT 81.020 119.390 81.190 119.560 ;
        RECT 81.020 119.030 81.190 119.200 ;
        RECT 81.020 118.670 81.190 118.840 ;
        RECT 81.020 118.310 81.190 118.480 ;
        RECT 81.020 117.950 81.190 118.120 ;
        RECT 81.020 117.590 81.190 117.760 ;
        RECT 81.570 120.245 81.740 120.415 ;
        RECT 81.570 119.885 81.740 120.055 ;
        RECT 81.570 119.525 81.740 119.695 ;
        RECT 81.570 119.165 81.740 119.335 ;
        RECT 81.570 118.805 81.740 118.975 ;
        RECT 81.570 118.445 81.740 118.615 ;
        RECT 81.570 118.085 81.740 118.255 ;
        RECT 81.570 117.725 81.740 117.895 ;
        RECT 82.740 120.245 82.910 120.415 ;
        RECT 82.740 119.885 82.910 120.055 ;
        RECT 82.740 119.525 82.910 119.695 ;
        RECT 82.740 119.165 82.910 119.335 ;
        RECT 82.740 118.805 82.910 118.975 ;
        RECT 84.310 120.370 84.480 120.540 ;
        RECT 84.310 120.010 84.480 120.180 ;
        RECT 84.310 119.650 84.480 119.820 ;
        RECT 84.310 119.290 84.480 119.460 ;
        RECT 84.310 118.930 84.480 119.100 ;
        RECT 85.480 120.370 85.650 120.540 ;
        RECT 85.480 120.010 85.650 120.180 ;
        RECT 85.480 119.650 85.650 119.820 ;
        RECT 85.480 119.290 85.650 119.460 ;
        RECT 85.480 118.930 85.650 119.100 ;
        RECT 86.030 120.470 86.200 120.640 ;
        RECT 86.030 120.110 86.200 120.280 ;
        RECT 86.030 119.750 86.200 119.920 ;
        RECT 86.030 119.390 86.200 119.560 ;
        RECT 86.030 119.030 86.200 119.200 ;
        RECT 82.740 118.445 82.910 118.615 ;
        RECT 84.895 118.510 85.065 118.680 ;
        RECT 86.030 118.670 86.200 118.840 ;
        RECT 86.030 118.310 86.200 118.480 ;
        RECT 82.740 118.085 82.910 118.255 ;
        RECT 82.740 117.725 82.910 117.895 ;
        RECT 84.310 118.090 84.480 118.260 ;
        RECT 84.310 117.730 84.480 117.900 ;
        RECT 81.020 117.230 81.190 117.400 ;
        RECT 82.155 117.350 82.325 117.520 ;
        RECT 84.310 117.370 84.480 117.540 ;
        RECT 81.020 116.870 81.190 117.040 ;
        RECT 81.020 116.510 81.190 116.680 ;
        RECT 81.020 116.150 81.190 116.320 ;
        RECT 81.020 115.790 81.190 115.960 ;
        RECT 81.020 115.430 81.190 115.600 ;
        RECT 81.020 115.070 81.190 115.240 ;
        RECT 81.020 114.710 81.190 114.880 ;
        RECT 81.020 114.350 81.190 114.520 ;
        RECT 81.570 116.965 81.740 117.135 ;
        RECT 81.570 116.605 81.740 116.775 ;
        RECT 81.570 116.245 81.740 116.415 ;
        RECT 81.570 115.885 81.740 116.055 ;
        RECT 81.570 115.525 81.740 115.695 ;
        RECT 81.570 115.165 81.740 115.335 ;
        RECT 81.570 114.805 81.740 114.975 ;
        RECT 81.570 114.445 81.740 114.615 ;
        RECT 82.740 116.965 82.910 117.135 ;
        RECT 82.740 116.605 82.910 116.775 ;
        RECT 84.310 117.010 84.480 117.180 ;
        RECT 84.310 116.650 84.480 116.820 ;
        RECT 85.480 118.090 85.650 118.260 ;
        RECT 85.480 117.730 85.650 117.900 ;
        RECT 85.480 117.370 85.650 117.540 ;
        RECT 85.480 117.010 85.650 117.180 ;
        RECT 85.480 116.650 85.650 116.820 ;
        RECT 86.030 117.950 86.200 118.120 ;
        RECT 86.030 117.590 86.200 117.760 ;
        RECT 87.960 138.290 88.130 138.460 ;
        RECT 88.320 138.290 88.490 138.460 ;
        RECT 88.680 138.290 88.850 138.460 ;
        RECT 89.040 138.290 89.210 138.460 ;
        RECT 89.400 138.290 89.570 138.460 ;
        RECT 89.760 138.290 89.930 138.460 ;
        RECT 90.120 138.290 90.290 138.460 ;
        RECT 87.660 137.940 87.830 138.110 ;
        RECT 90.430 137.940 90.600 138.110 ;
        RECT 87.660 137.580 87.830 137.750 ;
        RECT 88.865 137.620 89.035 137.790 ;
        RECT 89.225 137.620 89.395 137.790 ;
        RECT 90.430 137.580 90.600 137.750 ;
        RECT 87.660 137.220 87.830 137.390 ;
        RECT 87.660 136.860 87.830 137.030 ;
        RECT 87.660 136.500 87.830 136.670 ;
        RECT 87.660 136.140 87.830 136.310 ;
        RECT 87.660 135.780 87.830 135.950 ;
        RECT 87.660 135.420 87.830 135.590 ;
        RECT 88.210 137.235 88.380 137.405 ;
        RECT 88.210 136.875 88.380 137.045 ;
        RECT 88.210 136.515 88.380 136.685 ;
        RECT 89.880 137.235 90.050 137.405 ;
        RECT 89.880 136.875 90.050 137.045 ;
        RECT 89.880 136.515 90.050 136.685 ;
        RECT 88.865 136.340 89.035 136.510 ;
        RECT 89.225 136.340 89.395 136.510 ;
        RECT 88.210 136.155 88.380 136.325 ;
        RECT 88.210 135.795 88.380 135.965 ;
        RECT 88.210 135.435 88.380 135.605 ;
        RECT 89.880 136.155 90.050 136.325 ;
        RECT 89.880 135.795 90.050 135.965 ;
        RECT 89.880 135.435 90.050 135.605 ;
        RECT 90.430 137.220 90.600 137.390 ;
        RECT 90.430 136.860 90.600 137.030 ;
        RECT 90.430 136.500 90.600 136.670 ;
        RECT 90.430 136.140 90.600 136.310 ;
        RECT 90.430 135.780 90.600 135.950 ;
        RECT 90.430 135.420 90.600 135.590 ;
        RECT 87.660 135.060 87.830 135.230 ;
        RECT 88.865 135.060 89.035 135.230 ;
        RECT 89.225 135.060 89.395 135.230 ;
        RECT 90.430 135.060 90.600 135.230 ;
        RECT 87.660 134.700 87.830 134.870 ;
        RECT 87.660 134.340 87.830 134.510 ;
        RECT 87.660 133.980 87.830 134.150 ;
        RECT 87.660 133.620 87.830 133.790 ;
        RECT 87.660 133.260 87.830 133.430 ;
        RECT 88.210 134.640 88.380 134.810 ;
        RECT 88.210 134.280 88.380 134.450 ;
        RECT 88.210 133.920 88.380 134.090 ;
        RECT 88.210 133.560 88.380 133.730 ;
        RECT 88.210 133.200 88.380 133.370 ;
        RECT 89.880 134.640 90.050 134.810 ;
        RECT 89.880 134.280 90.050 134.450 ;
        RECT 89.880 133.920 90.050 134.090 ;
        RECT 89.880 133.560 90.050 133.730 ;
        RECT 89.880 133.200 90.050 133.370 ;
        RECT 90.430 134.700 90.600 134.870 ;
        RECT 90.430 134.340 90.600 134.510 ;
        RECT 90.430 133.980 90.600 134.150 ;
        RECT 90.430 133.620 90.600 133.790 ;
        RECT 90.430 133.260 90.600 133.430 ;
        RECT 87.660 132.900 87.830 133.070 ;
        RECT 88.865 132.780 89.035 132.950 ;
        RECT 89.225 132.780 89.395 132.950 ;
        RECT 90.430 132.900 90.600 133.070 ;
        RECT 87.660 132.540 87.830 132.710 ;
        RECT 90.430 132.540 90.600 132.710 ;
        RECT 87.660 132.180 87.830 132.350 ;
        RECT 87.660 131.820 87.830 131.990 ;
        RECT 87.660 131.460 87.830 131.630 ;
        RECT 87.660 131.100 87.830 131.270 ;
        RECT 88.210 132.360 88.380 132.530 ;
        RECT 88.210 132.000 88.380 132.170 ;
        RECT 88.210 131.640 88.380 131.810 ;
        RECT 88.210 131.280 88.380 131.450 ;
        RECT 88.210 130.920 88.380 131.090 ;
        RECT 89.880 132.360 90.050 132.530 ;
        RECT 89.880 132.000 90.050 132.170 ;
        RECT 89.880 131.640 90.050 131.810 ;
        RECT 89.880 131.280 90.050 131.450 ;
        RECT 89.880 130.920 90.050 131.090 ;
        RECT 90.430 132.180 90.600 132.350 ;
        RECT 90.430 131.820 90.600 131.990 ;
        RECT 90.430 131.460 90.600 131.630 ;
        RECT 90.430 131.100 90.600 131.270 ;
        RECT 87.660 130.740 87.830 130.910 ;
        RECT 90.430 130.740 90.600 130.910 ;
        RECT 87.660 130.380 87.830 130.550 ;
        RECT 88.865 130.500 89.035 130.670 ;
        RECT 89.225 130.500 89.395 130.670 ;
        RECT 90.430 130.380 90.600 130.550 ;
        RECT 87.660 130.020 87.830 130.190 ;
        RECT 87.660 129.660 87.830 129.830 ;
        RECT 87.660 129.300 87.830 129.470 ;
        RECT 87.660 128.940 87.830 129.110 ;
        RECT 87.660 128.580 87.830 128.750 ;
        RECT 87.660 128.220 87.830 128.390 ;
        RECT 88.210 130.115 88.380 130.285 ;
        RECT 88.210 129.755 88.380 129.925 ;
        RECT 88.210 129.395 88.380 129.565 ;
        RECT 89.880 130.115 90.050 130.285 ;
        RECT 89.880 129.755 90.050 129.925 ;
        RECT 89.880 129.395 90.050 129.565 ;
        RECT 88.865 129.220 89.035 129.390 ;
        RECT 89.225 129.220 89.395 129.390 ;
        RECT 88.210 129.035 88.380 129.205 ;
        RECT 88.210 128.675 88.380 128.845 ;
        RECT 88.210 128.315 88.380 128.485 ;
        RECT 89.880 129.035 90.050 129.205 ;
        RECT 89.880 128.675 90.050 128.845 ;
        RECT 89.880 128.315 90.050 128.485 ;
        RECT 90.430 130.020 90.600 130.190 ;
        RECT 90.430 129.660 90.600 129.830 ;
        RECT 90.430 129.300 90.600 129.470 ;
        RECT 90.430 128.940 90.600 129.110 ;
        RECT 90.430 128.580 90.600 128.750 ;
        RECT 90.430 128.220 90.600 128.390 ;
        RECT 87.660 127.860 87.830 128.030 ;
        RECT 88.865 127.940 89.035 128.110 ;
        RECT 89.225 127.940 89.395 128.110 ;
        RECT 90.430 127.860 90.600 128.030 ;
        RECT 87.660 127.500 87.830 127.670 ;
        RECT 87.660 127.140 87.830 127.310 ;
        RECT 87.660 126.780 87.830 126.950 ;
        RECT 87.660 126.420 87.830 126.590 ;
        RECT 87.660 126.060 87.830 126.230 ;
        RECT 87.660 125.700 87.830 125.870 ;
        RECT 88.210 127.555 88.380 127.725 ;
        RECT 88.210 127.195 88.380 127.365 ;
        RECT 88.210 126.835 88.380 127.005 ;
        RECT 89.880 127.555 90.050 127.725 ;
        RECT 89.880 127.195 90.050 127.365 ;
        RECT 89.880 126.835 90.050 127.005 ;
        RECT 88.865 126.660 89.035 126.830 ;
        RECT 89.225 126.660 89.395 126.830 ;
        RECT 88.210 126.475 88.380 126.645 ;
        RECT 88.210 126.115 88.380 126.285 ;
        RECT 88.210 125.755 88.380 125.925 ;
        RECT 89.880 126.475 90.050 126.645 ;
        RECT 89.880 126.115 90.050 126.285 ;
        RECT 89.880 125.755 90.050 125.925 ;
        RECT 90.430 127.500 90.600 127.670 ;
        RECT 90.430 127.140 90.600 127.310 ;
        RECT 90.430 126.780 90.600 126.950 ;
        RECT 90.430 126.420 90.600 126.590 ;
        RECT 90.430 126.060 90.600 126.230 ;
        RECT 90.430 125.700 90.600 125.870 ;
        RECT 87.660 125.340 87.830 125.510 ;
        RECT 88.865 125.380 89.035 125.550 ;
        RECT 89.225 125.380 89.395 125.550 ;
        RECT 87.660 124.980 87.830 125.150 ;
        RECT 90.430 125.340 90.600 125.510 ;
        RECT 87.660 124.620 87.830 124.790 ;
        RECT 87.660 124.260 87.830 124.430 ;
        RECT 87.660 123.900 87.830 124.070 ;
        RECT 87.660 123.540 87.830 123.710 ;
        RECT 88.210 124.960 88.380 125.130 ;
        RECT 88.210 124.600 88.380 124.770 ;
        RECT 88.210 124.240 88.380 124.410 ;
        RECT 88.210 123.880 88.380 124.050 ;
        RECT 88.210 123.520 88.380 123.690 ;
        RECT 90.430 124.980 90.600 125.150 ;
        RECT 90.430 124.620 90.600 124.790 ;
        RECT 90.430 124.260 90.600 124.430 ;
        RECT 90.430 123.900 90.600 124.070 ;
        RECT 90.430 123.540 90.600 123.710 ;
        RECT 87.660 123.180 87.830 123.350 ;
        RECT 88.865 123.100 89.035 123.270 ;
        RECT 89.225 123.100 89.395 123.270 ;
        RECT 90.430 123.180 90.600 123.350 ;
        RECT 87.660 122.820 87.830 122.990 ;
        RECT 87.660 122.460 87.830 122.630 ;
        RECT 87.660 122.100 87.830 122.270 ;
        RECT 87.660 121.740 87.830 121.910 ;
        RECT 87.660 121.380 87.830 121.550 ;
        RECT 88.210 122.680 88.380 122.850 ;
        RECT 88.210 122.320 88.380 122.490 ;
        RECT 88.210 121.960 88.380 122.130 ;
        RECT 88.210 121.600 88.380 121.770 ;
        RECT 88.210 121.240 88.380 121.410 ;
        RECT 90.430 122.820 90.600 122.990 ;
        RECT 90.430 122.460 90.600 122.630 ;
        RECT 90.430 122.100 90.600 122.270 ;
        RECT 90.430 121.740 90.600 121.910 ;
        RECT 90.430 121.380 90.600 121.550 ;
        RECT 87.660 121.020 87.830 121.190 ;
        RECT 90.430 121.020 90.600 121.190 ;
        RECT 87.660 120.660 87.830 120.830 ;
        RECT 88.865 120.820 89.035 120.990 ;
        RECT 89.225 120.820 89.395 120.990 ;
        RECT 90.430 120.660 90.600 120.830 ;
        RECT 87.660 120.300 87.830 120.470 ;
        RECT 87.660 119.940 87.830 120.110 ;
        RECT 87.660 119.580 87.830 119.750 ;
        RECT 87.660 119.220 87.830 119.390 ;
        RECT 87.660 118.860 87.830 119.030 ;
        RECT 87.660 118.500 87.830 118.670 ;
        RECT 88.210 120.435 88.380 120.605 ;
        RECT 88.210 120.075 88.380 120.245 ;
        RECT 88.210 119.715 88.380 119.885 ;
        RECT 89.880 120.435 90.050 120.605 ;
        RECT 89.880 120.075 90.050 120.245 ;
        RECT 89.880 119.715 90.050 119.885 ;
        RECT 88.865 119.540 89.035 119.710 ;
        RECT 89.225 119.540 89.395 119.710 ;
        RECT 88.210 119.355 88.380 119.525 ;
        RECT 88.210 118.995 88.380 119.165 ;
        RECT 88.210 118.635 88.380 118.805 ;
        RECT 89.880 119.355 90.050 119.525 ;
        RECT 89.880 118.995 90.050 119.165 ;
        RECT 89.880 118.635 90.050 118.805 ;
        RECT 90.430 120.300 90.600 120.470 ;
        RECT 90.430 119.940 90.600 120.110 ;
        RECT 90.430 119.580 90.600 119.750 ;
        RECT 90.430 119.220 90.600 119.390 ;
        RECT 90.430 118.860 90.600 119.030 ;
        RECT 90.430 118.500 90.600 118.670 ;
        RECT 87.660 118.140 87.830 118.310 ;
        RECT 88.865 118.260 89.035 118.430 ;
        RECT 89.225 118.260 89.395 118.430 ;
        RECT 90.430 118.140 90.600 118.310 ;
        RECT 87.960 117.590 88.130 117.760 ;
        RECT 88.320 117.590 88.490 117.760 ;
        RECT 88.680 117.590 88.850 117.760 ;
        RECT 89.040 117.590 89.210 117.760 ;
        RECT 89.400 117.590 89.570 117.760 ;
        RECT 89.760 117.590 89.930 117.760 ;
        RECT 90.120 117.590 90.290 117.760 ;
        RECT 92.215 138.290 92.385 138.460 ;
        RECT 92.575 138.290 92.745 138.460 ;
        RECT 92.935 138.290 93.105 138.460 ;
        RECT 93.295 138.290 93.465 138.460 ;
        RECT 93.655 138.290 93.825 138.460 ;
        RECT 91.915 137.940 92.085 138.110 ;
        RECT 94.185 137.940 94.355 138.110 ;
        RECT 91.915 137.580 92.085 137.750 ;
        RECT 93.050 137.620 93.220 137.790 ;
        RECT 94.185 137.580 94.355 137.750 ;
        RECT 91.915 137.220 92.085 137.390 ;
        RECT 91.915 136.860 92.085 137.030 ;
        RECT 91.915 136.500 92.085 136.670 ;
        RECT 91.915 136.140 92.085 136.310 ;
        RECT 91.915 135.780 92.085 135.950 ;
        RECT 91.915 135.420 92.085 135.590 ;
        RECT 92.465 137.235 92.635 137.405 ;
        RECT 92.465 136.875 92.635 137.045 ;
        RECT 92.465 136.515 92.635 136.685 ;
        RECT 93.635 137.235 93.805 137.405 ;
        RECT 93.635 136.875 93.805 137.045 ;
        RECT 93.635 136.515 93.805 136.685 ;
        RECT 93.050 136.340 93.220 136.510 ;
        RECT 92.465 136.155 92.635 136.325 ;
        RECT 92.465 135.795 92.635 135.965 ;
        RECT 92.465 135.435 92.635 135.605 ;
        RECT 93.635 136.155 93.805 136.325 ;
        RECT 93.635 135.795 93.805 135.965 ;
        RECT 93.635 135.435 93.805 135.605 ;
        RECT 94.185 137.220 94.355 137.390 ;
        RECT 94.185 136.860 94.355 137.030 ;
        RECT 94.185 136.500 94.355 136.670 ;
        RECT 94.185 136.140 94.355 136.310 ;
        RECT 94.185 135.780 94.355 135.950 ;
        RECT 94.185 135.420 94.355 135.590 ;
        RECT 91.915 135.060 92.085 135.230 ;
        RECT 93.050 135.060 93.220 135.230 ;
        RECT 94.185 135.060 94.355 135.230 ;
        RECT 91.915 134.700 92.085 134.870 ;
        RECT 91.915 134.340 92.085 134.510 ;
        RECT 91.915 133.980 92.085 134.150 ;
        RECT 91.915 133.620 92.085 133.790 ;
        RECT 91.915 133.260 92.085 133.430 ;
        RECT 92.465 134.640 92.635 134.810 ;
        RECT 92.465 134.280 92.635 134.450 ;
        RECT 92.465 133.920 92.635 134.090 ;
        RECT 92.465 133.560 92.635 133.730 ;
        RECT 92.465 133.200 92.635 133.370 ;
        RECT 93.635 134.640 93.805 134.810 ;
        RECT 93.635 134.280 93.805 134.450 ;
        RECT 93.635 133.920 93.805 134.090 ;
        RECT 93.635 133.560 93.805 133.730 ;
        RECT 93.635 133.200 93.805 133.370 ;
        RECT 94.185 134.700 94.355 134.870 ;
        RECT 94.185 134.340 94.355 134.510 ;
        RECT 94.185 133.980 94.355 134.150 ;
        RECT 94.185 133.620 94.355 133.790 ;
        RECT 94.185 133.260 94.355 133.430 ;
        RECT 91.915 132.900 92.085 133.070 ;
        RECT 93.050 132.780 93.220 132.950 ;
        RECT 94.185 132.900 94.355 133.070 ;
        RECT 91.915 132.540 92.085 132.710 ;
        RECT 94.185 132.540 94.355 132.710 ;
        RECT 91.915 132.180 92.085 132.350 ;
        RECT 91.915 131.820 92.085 131.990 ;
        RECT 91.915 131.460 92.085 131.630 ;
        RECT 91.915 131.100 92.085 131.270 ;
        RECT 92.465 132.360 92.635 132.530 ;
        RECT 92.465 132.000 92.635 132.170 ;
        RECT 92.465 131.640 92.635 131.810 ;
        RECT 92.465 131.280 92.635 131.450 ;
        RECT 92.465 130.920 92.635 131.090 ;
        RECT 93.635 132.360 93.805 132.530 ;
        RECT 93.635 132.000 93.805 132.170 ;
        RECT 93.635 131.640 93.805 131.810 ;
        RECT 93.635 131.280 93.805 131.450 ;
        RECT 93.635 130.920 93.805 131.090 ;
        RECT 94.185 132.180 94.355 132.350 ;
        RECT 94.185 131.820 94.355 131.990 ;
        RECT 94.185 131.460 94.355 131.630 ;
        RECT 94.185 131.100 94.355 131.270 ;
        RECT 91.915 130.740 92.085 130.910 ;
        RECT 94.185 130.740 94.355 130.910 ;
        RECT 91.915 130.380 92.085 130.550 ;
        RECT 93.050 130.500 93.220 130.670 ;
        RECT 94.185 130.380 94.355 130.550 ;
        RECT 91.915 130.020 92.085 130.190 ;
        RECT 91.915 129.660 92.085 129.830 ;
        RECT 91.915 129.300 92.085 129.470 ;
        RECT 91.915 128.940 92.085 129.110 ;
        RECT 91.915 128.580 92.085 128.750 ;
        RECT 91.915 128.220 92.085 128.390 ;
        RECT 92.465 130.115 92.635 130.285 ;
        RECT 92.465 129.755 92.635 129.925 ;
        RECT 92.465 129.395 92.635 129.565 ;
        RECT 93.635 130.115 93.805 130.285 ;
        RECT 93.635 129.755 93.805 129.925 ;
        RECT 93.635 129.395 93.805 129.565 ;
        RECT 93.050 129.220 93.220 129.390 ;
        RECT 92.465 129.035 92.635 129.205 ;
        RECT 92.465 128.675 92.635 128.845 ;
        RECT 92.465 128.315 92.635 128.485 ;
        RECT 93.635 129.035 93.805 129.205 ;
        RECT 93.635 128.675 93.805 128.845 ;
        RECT 93.635 128.315 93.805 128.485 ;
        RECT 94.185 130.020 94.355 130.190 ;
        RECT 94.185 129.660 94.355 129.830 ;
        RECT 94.185 129.300 94.355 129.470 ;
        RECT 94.185 128.940 94.355 129.110 ;
        RECT 94.185 128.580 94.355 128.750 ;
        RECT 94.185 128.220 94.355 128.390 ;
        RECT 91.915 127.860 92.085 128.030 ;
        RECT 93.050 127.940 93.220 128.110 ;
        RECT 94.185 127.860 94.355 128.030 ;
        RECT 91.915 127.500 92.085 127.670 ;
        RECT 91.915 127.140 92.085 127.310 ;
        RECT 91.915 126.780 92.085 126.950 ;
        RECT 91.915 126.420 92.085 126.590 ;
        RECT 91.915 126.060 92.085 126.230 ;
        RECT 91.915 125.700 92.085 125.870 ;
        RECT 92.465 127.555 92.635 127.725 ;
        RECT 92.465 127.195 92.635 127.365 ;
        RECT 92.465 126.835 92.635 127.005 ;
        RECT 93.635 127.555 93.805 127.725 ;
        RECT 93.635 127.195 93.805 127.365 ;
        RECT 93.635 126.835 93.805 127.005 ;
        RECT 93.050 126.660 93.220 126.830 ;
        RECT 92.465 126.475 92.635 126.645 ;
        RECT 92.465 126.115 92.635 126.285 ;
        RECT 92.465 125.755 92.635 125.925 ;
        RECT 93.635 126.475 93.805 126.645 ;
        RECT 93.635 126.115 93.805 126.285 ;
        RECT 93.635 125.755 93.805 125.925 ;
        RECT 94.185 127.500 94.355 127.670 ;
        RECT 94.185 127.140 94.355 127.310 ;
        RECT 94.185 126.780 94.355 126.950 ;
        RECT 94.185 126.420 94.355 126.590 ;
        RECT 94.185 126.060 94.355 126.230 ;
        RECT 94.185 125.700 94.355 125.870 ;
        RECT 91.915 125.340 92.085 125.510 ;
        RECT 93.050 125.380 93.220 125.550 ;
        RECT 91.915 124.980 92.085 125.150 ;
        RECT 94.185 125.340 94.355 125.510 ;
        RECT 91.915 124.620 92.085 124.790 ;
        RECT 91.915 124.260 92.085 124.430 ;
        RECT 91.915 123.900 92.085 124.070 ;
        RECT 91.915 123.540 92.085 123.710 ;
        RECT 93.635 124.960 93.805 125.130 ;
        RECT 93.635 124.600 93.805 124.770 ;
        RECT 93.635 124.240 93.805 124.410 ;
        RECT 93.635 123.880 93.805 124.050 ;
        RECT 93.635 123.520 93.805 123.690 ;
        RECT 94.185 124.980 94.355 125.150 ;
        RECT 94.185 124.620 94.355 124.790 ;
        RECT 94.185 124.260 94.355 124.430 ;
        RECT 94.185 123.900 94.355 124.070 ;
        RECT 94.185 123.540 94.355 123.710 ;
        RECT 91.915 123.180 92.085 123.350 ;
        RECT 93.050 123.100 93.220 123.270 ;
        RECT 94.185 123.180 94.355 123.350 ;
        RECT 91.915 122.820 92.085 122.990 ;
        RECT 91.915 122.460 92.085 122.630 ;
        RECT 91.915 122.100 92.085 122.270 ;
        RECT 91.915 121.740 92.085 121.910 ;
        RECT 91.915 121.380 92.085 121.550 ;
        RECT 93.635 122.680 93.805 122.850 ;
        RECT 93.635 122.320 93.805 122.490 ;
        RECT 93.635 121.960 93.805 122.130 ;
        RECT 93.635 121.600 93.805 121.770 ;
        RECT 93.635 121.240 93.805 121.410 ;
        RECT 94.185 122.820 94.355 122.990 ;
        RECT 94.185 122.460 94.355 122.630 ;
        RECT 94.185 122.100 94.355 122.270 ;
        RECT 94.185 121.740 94.355 121.910 ;
        RECT 94.185 121.380 94.355 121.550 ;
        RECT 91.915 121.020 92.085 121.190 ;
        RECT 94.185 121.020 94.355 121.190 ;
        RECT 91.915 120.660 92.085 120.830 ;
        RECT 93.050 120.820 93.220 120.990 ;
        RECT 94.185 120.660 94.355 120.830 ;
        RECT 91.915 120.300 92.085 120.470 ;
        RECT 91.915 119.940 92.085 120.110 ;
        RECT 91.915 119.580 92.085 119.750 ;
        RECT 91.915 119.220 92.085 119.390 ;
        RECT 91.915 118.860 92.085 119.030 ;
        RECT 91.915 118.500 92.085 118.670 ;
        RECT 92.465 120.435 92.635 120.605 ;
        RECT 92.465 120.075 92.635 120.245 ;
        RECT 92.465 119.715 92.635 119.885 ;
        RECT 93.635 120.435 93.805 120.605 ;
        RECT 93.635 120.075 93.805 120.245 ;
        RECT 93.635 119.715 93.805 119.885 ;
        RECT 93.050 119.540 93.220 119.710 ;
        RECT 92.465 119.355 92.635 119.525 ;
        RECT 92.465 118.995 92.635 119.165 ;
        RECT 92.465 118.635 92.635 118.805 ;
        RECT 93.635 119.355 93.805 119.525 ;
        RECT 93.635 118.995 93.805 119.165 ;
        RECT 93.635 118.635 93.805 118.805 ;
        RECT 94.185 120.300 94.355 120.470 ;
        RECT 94.185 119.940 94.355 120.110 ;
        RECT 94.185 119.580 94.355 119.750 ;
        RECT 94.185 119.220 94.355 119.390 ;
        RECT 94.185 118.860 94.355 119.030 ;
        RECT 94.185 118.500 94.355 118.670 ;
        RECT 91.915 118.140 92.085 118.310 ;
        RECT 93.050 118.260 93.220 118.430 ;
        RECT 94.185 118.140 94.355 118.310 ;
        RECT 92.215 117.590 92.385 117.760 ;
        RECT 92.575 117.590 92.745 117.760 ;
        RECT 92.935 117.590 93.105 117.760 ;
        RECT 93.295 117.590 93.465 117.760 ;
        RECT 93.655 117.590 93.825 117.760 ;
        RECT 96.080 138.190 96.250 138.360 ;
        RECT 96.080 137.830 96.250 138.000 ;
        RECT 96.080 137.470 96.250 137.640 ;
        RECT 96.630 138.890 96.800 139.060 ;
        RECT 96.630 138.530 96.800 138.700 ;
        RECT 96.630 138.170 96.800 138.340 ;
        RECT 96.630 137.810 96.800 137.980 ;
        RECT 96.630 137.450 96.800 137.620 ;
        RECT 98.300 138.890 98.470 139.060 ;
        RECT 98.300 138.530 98.470 138.700 ;
        RECT 98.300 138.170 98.470 138.340 ;
        RECT 98.300 137.810 98.470 137.980 ;
        RECT 98.300 137.450 98.470 137.620 ;
        RECT 100.220 138.890 100.390 139.060 ;
        RECT 100.220 138.530 100.390 138.700 ;
        RECT 100.220 138.170 100.390 138.340 ;
        RECT 100.220 137.810 100.390 137.980 ;
        RECT 100.220 137.450 100.390 137.620 ;
        RECT 102.440 138.910 102.610 139.080 ;
        RECT 102.440 138.550 102.610 138.720 ;
        RECT 102.440 138.190 102.610 138.360 ;
        RECT 102.440 137.830 102.610 138.000 ;
        RECT 102.440 137.470 102.610 137.640 ;
        RECT 96.080 137.110 96.250 137.280 ;
        RECT 97.285 137.030 97.455 137.200 ;
        RECT 97.645 137.030 97.815 137.200 ;
        RECT 100.875 137.030 101.045 137.200 ;
        RECT 101.235 137.030 101.405 137.200 ;
        RECT 102.440 137.110 102.610 137.280 ;
        RECT 96.080 136.750 96.250 136.920 ;
        RECT 96.080 136.390 96.250 136.560 ;
        RECT 96.080 136.030 96.250 136.200 ;
        RECT 96.080 135.670 96.250 135.840 ;
        RECT 96.080 135.310 96.250 135.480 ;
        RECT 96.630 136.610 96.800 136.780 ;
        RECT 96.630 136.250 96.800 136.420 ;
        RECT 96.630 135.890 96.800 136.060 ;
        RECT 96.630 135.530 96.800 135.700 ;
        RECT 96.630 135.170 96.800 135.340 ;
        RECT 98.300 136.610 98.470 136.780 ;
        RECT 98.300 136.250 98.470 136.420 ;
        RECT 98.300 135.890 98.470 136.060 ;
        RECT 98.300 135.530 98.470 135.700 ;
        RECT 98.300 135.170 98.470 135.340 ;
        RECT 100.220 136.610 100.390 136.780 ;
        RECT 100.220 136.250 100.390 136.420 ;
        RECT 100.220 135.890 100.390 136.060 ;
        RECT 100.220 135.530 100.390 135.700 ;
        RECT 100.220 135.170 100.390 135.340 ;
        RECT 102.440 136.750 102.610 136.920 ;
        RECT 102.440 136.390 102.610 136.560 ;
        RECT 102.440 136.030 102.610 136.200 ;
        RECT 102.440 135.670 102.610 135.840 ;
        RECT 102.440 135.310 102.610 135.480 ;
        RECT 96.080 134.950 96.250 135.120 ;
        RECT 102.440 134.950 102.610 135.120 ;
        RECT 96.080 134.590 96.250 134.760 ;
        RECT 97.285 134.750 97.455 134.920 ;
        RECT 97.645 134.750 97.815 134.920 ;
        RECT 100.875 134.750 101.045 134.920 ;
        RECT 101.235 134.750 101.405 134.920 ;
        RECT 102.440 134.590 102.610 134.760 ;
        RECT 96.080 134.230 96.250 134.400 ;
        RECT 96.080 133.870 96.250 134.040 ;
        RECT 96.080 133.510 96.250 133.680 ;
        RECT 96.080 133.150 96.250 133.320 ;
        RECT 96.080 132.790 96.250 132.960 ;
        RECT 96.630 134.330 96.800 134.500 ;
        RECT 96.630 133.970 96.800 134.140 ;
        RECT 96.630 133.610 96.800 133.780 ;
        RECT 96.630 133.250 96.800 133.420 ;
        RECT 96.630 132.890 96.800 133.060 ;
        RECT 98.300 134.330 98.470 134.500 ;
        RECT 98.300 133.970 98.470 134.140 ;
        RECT 98.300 133.610 98.470 133.780 ;
        RECT 98.300 133.250 98.470 133.420 ;
        RECT 98.300 132.890 98.470 133.060 ;
        RECT 100.220 134.330 100.390 134.500 ;
        RECT 100.220 133.970 100.390 134.140 ;
        RECT 100.220 133.610 100.390 133.780 ;
        RECT 100.220 133.250 100.390 133.420 ;
        RECT 100.220 132.890 100.390 133.060 ;
        RECT 102.440 134.230 102.610 134.400 ;
        RECT 102.440 133.870 102.610 134.040 ;
        RECT 102.440 133.510 102.610 133.680 ;
        RECT 102.440 133.150 102.610 133.320 ;
        RECT 102.440 132.790 102.610 132.960 ;
        RECT 96.080 132.430 96.250 132.600 ;
        RECT 97.285 132.470 97.455 132.640 ;
        RECT 97.645 132.470 97.815 132.640 ;
        RECT 100.875 132.470 101.045 132.640 ;
        RECT 101.235 132.470 101.405 132.640 ;
        RECT 96.080 132.070 96.250 132.240 ;
        RECT 102.440 132.430 102.610 132.600 ;
        RECT 96.080 131.710 96.250 131.880 ;
        RECT 96.080 131.350 96.250 131.520 ;
        RECT 96.080 130.990 96.250 131.160 ;
        RECT 96.080 130.630 96.250 130.800 ;
        RECT 96.630 132.050 96.800 132.220 ;
        RECT 96.630 131.690 96.800 131.860 ;
        RECT 96.630 131.330 96.800 131.500 ;
        RECT 96.630 130.970 96.800 131.140 ;
        RECT 96.630 130.610 96.800 130.780 ;
        RECT 98.300 132.050 98.470 132.220 ;
        RECT 98.300 131.690 98.470 131.860 ;
        RECT 98.300 131.330 98.470 131.500 ;
        RECT 98.300 130.970 98.470 131.140 ;
        RECT 98.300 130.610 98.470 130.780 ;
        RECT 100.220 132.050 100.390 132.220 ;
        RECT 100.220 131.690 100.390 131.860 ;
        RECT 100.220 131.330 100.390 131.500 ;
        RECT 100.220 130.970 100.390 131.140 ;
        RECT 100.220 130.610 100.390 130.780 ;
        RECT 102.440 132.070 102.610 132.240 ;
        RECT 102.440 131.710 102.610 131.880 ;
        RECT 102.440 131.350 102.610 131.520 ;
        RECT 102.440 130.990 102.610 131.160 ;
        RECT 102.440 130.630 102.610 130.800 ;
        RECT 96.080 130.270 96.250 130.440 ;
        RECT 97.285 130.190 97.455 130.360 ;
        RECT 97.645 130.190 97.815 130.360 ;
        RECT 100.875 130.190 101.045 130.360 ;
        RECT 101.235 130.190 101.405 130.360 ;
        RECT 102.440 130.270 102.610 130.440 ;
        RECT 96.080 129.910 96.250 130.080 ;
        RECT 96.080 129.550 96.250 129.720 ;
        RECT 96.080 129.190 96.250 129.360 ;
        RECT 96.080 128.830 96.250 129.000 ;
        RECT 96.080 128.470 96.250 128.640 ;
        RECT 96.630 129.770 96.800 129.940 ;
        RECT 96.630 129.410 96.800 129.580 ;
        RECT 96.630 129.050 96.800 129.220 ;
        RECT 96.630 128.690 96.800 128.860 ;
        RECT 96.630 128.330 96.800 128.500 ;
        RECT 98.300 129.770 98.470 129.940 ;
        RECT 98.300 129.410 98.470 129.580 ;
        RECT 98.300 129.050 98.470 129.220 ;
        RECT 98.300 128.690 98.470 128.860 ;
        RECT 98.300 128.330 98.470 128.500 ;
        RECT 101.890 129.770 102.060 129.940 ;
        RECT 101.890 129.410 102.060 129.580 ;
        RECT 101.890 129.050 102.060 129.220 ;
        RECT 101.890 128.690 102.060 128.860 ;
        RECT 101.890 128.330 102.060 128.500 ;
        RECT 102.440 129.910 102.610 130.080 ;
        RECT 102.440 129.550 102.610 129.720 ;
        RECT 102.440 129.190 102.610 129.360 ;
        RECT 102.440 128.830 102.610 129.000 ;
        RECT 102.440 128.470 102.610 128.640 ;
        RECT 96.080 128.110 96.250 128.280 ;
        RECT 102.440 128.110 102.610 128.280 ;
        RECT 96.080 127.750 96.250 127.920 ;
        RECT 97.285 127.910 97.455 128.080 ;
        RECT 97.645 127.910 97.815 128.080 ;
        RECT 100.875 127.910 101.045 128.080 ;
        RECT 101.235 127.910 101.405 128.080 ;
        RECT 102.440 127.750 102.610 127.920 ;
        RECT 96.080 127.390 96.250 127.560 ;
        RECT 96.080 127.030 96.250 127.200 ;
        RECT 96.080 126.670 96.250 126.840 ;
        RECT 96.080 126.310 96.250 126.480 ;
        RECT 96.080 125.950 96.250 126.120 ;
        RECT 96.630 127.490 96.800 127.660 ;
        RECT 96.630 127.130 96.800 127.300 ;
        RECT 96.630 126.770 96.800 126.940 ;
        RECT 96.630 126.410 96.800 126.580 ;
        RECT 96.630 126.050 96.800 126.220 ;
        RECT 98.300 127.490 98.470 127.660 ;
        RECT 98.300 127.130 98.470 127.300 ;
        RECT 98.300 126.770 98.470 126.940 ;
        RECT 98.300 126.410 98.470 126.580 ;
        RECT 98.300 126.050 98.470 126.220 ;
        RECT 101.890 127.490 102.060 127.660 ;
        RECT 101.890 127.130 102.060 127.300 ;
        RECT 101.890 126.770 102.060 126.940 ;
        RECT 101.890 126.410 102.060 126.580 ;
        RECT 101.890 126.050 102.060 126.220 ;
        RECT 102.440 127.390 102.610 127.560 ;
        RECT 102.440 127.030 102.610 127.200 ;
        RECT 102.440 126.670 102.610 126.840 ;
        RECT 102.440 126.310 102.610 126.480 ;
        RECT 102.440 125.950 102.610 126.120 ;
        RECT 96.080 125.590 96.250 125.760 ;
        RECT 97.285 125.630 97.455 125.800 ;
        RECT 97.645 125.630 97.815 125.800 ;
        RECT 100.875 125.630 101.045 125.800 ;
        RECT 101.235 125.630 101.405 125.800 ;
        RECT 96.080 125.230 96.250 125.400 ;
        RECT 102.440 125.590 102.610 125.760 ;
        RECT 96.080 124.870 96.250 125.040 ;
        RECT 96.080 124.510 96.250 124.680 ;
        RECT 96.080 124.150 96.250 124.320 ;
        RECT 96.080 123.790 96.250 123.960 ;
        RECT 96.630 125.210 96.800 125.380 ;
        RECT 96.630 124.850 96.800 125.020 ;
        RECT 96.630 124.490 96.800 124.660 ;
        RECT 96.630 124.130 96.800 124.300 ;
        RECT 96.630 123.770 96.800 123.940 ;
        RECT 98.300 125.210 98.470 125.380 ;
        RECT 98.300 124.850 98.470 125.020 ;
        RECT 98.300 124.490 98.470 124.660 ;
        RECT 98.300 124.130 98.470 124.300 ;
        RECT 98.300 123.770 98.470 123.940 ;
        RECT 100.220 125.210 100.390 125.380 ;
        RECT 100.220 124.850 100.390 125.020 ;
        RECT 100.220 124.490 100.390 124.660 ;
        RECT 100.220 124.130 100.390 124.300 ;
        RECT 100.220 123.770 100.390 123.940 ;
        RECT 102.440 125.230 102.610 125.400 ;
        RECT 102.440 124.870 102.610 125.040 ;
        RECT 102.440 124.510 102.610 124.680 ;
        RECT 102.440 124.150 102.610 124.320 ;
        RECT 102.440 123.790 102.610 123.960 ;
        RECT 96.080 123.430 96.250 123.600 ;
        RECT 97.285 123.350 97.455 123.520 ;
        RECT 97.645 123.350 97.815 123.520 ;
        RECT 100.875 123.350 101.045 123.520 ;
        RECT 101.235 123.350 101.405 123.520 ;
        RECT 102.440 123.430 102.610 123.600 ;
        RECT 96.080 123.070 96.250 123.240 ;
        RECT 96.080 122.710 96.250 122.880 ;
        RECT 96.080 122.350 96.250 122.520 ;
        RECT 96.080 121.990 96.250 122.160 ;
        RECT 96.080 121.630 96.250 121.800 ;
        RECT 96.630 122.930 96.800 123.100 ;
        RECT 96.630 122.570 96.800 122.740 ;
        RECT 96.630 122.210 96.800 122.380 ;
        RECT 96.630 121.850 96.800 122.020 ;
        RECT 96.630 121.490 96.800 121.660 ;
        RECT 98.300 122.930 98.470 123.100 ;
        RECT 98.300 122.570 98.470 122.740 ;
        RECT 98.300 122.210 98.470 122.380 ;
        RECT 98.300 121.850 98.470 122.020 ;
        RECT 98.300 121.490 98.470 121.660 ;
        RECT 100.220 122.930 100.390 123.100 ;
        RECT 100.220 122.570 100.390 122.740 ;
        RECT 100.220 122.210 100.390 122.380 ;
        RECT 100.220 121.850 100.390 122.020 ;
        RECT 100.220 121.490 100.390 121.660 ;
        RECT 102.440 123.070 102.610 123.240 ;
        RECT 102.440 122.710 102.610 122.880 ;
        RECT 102.440 122.350 102.610 122.520 ;
        RECT 102.440 121.990 102.610 122.160 ;
        RECT 102.440 121.630 102.610 121.800 ;
        RECT 96.080 121.270 96.250 121.440 ;
        RECT 102.440 121.270 102.610 121.440 ;
        RECT 96.080 120.910 96.250 121.080 ;
        RECT 97.285 121.070 97.455 121.240 ;
        RECT 97.645 121.070 97.815 121.240 ;
        RECT 100.875 121.070 101.045 121.240 ;
        RECT 101.235 121.070 101.405 121.240 ;
        RECT 102.440 120.910 102.610 121.080 ;
        RECT 96.080 120.550 96.250 120.720 ;
        RECT 96.080 120.190 96.250 120.360 ;
        RECT 96.080 119.830 96.250 120.000 ;
        RECT 96.080 119.470 96.250 119.640 ;
        RECT 96.080 119.110 96.250 119.280 ;
        RECT 96.630 120.650 96.800 120.820 ;
        RECT 96.630 120.290 96.800 120.460 ;
        RECT 96.630 119.930 96.800 120.100 ;
        RECT 96.630 119.570 96.800 119.740 ;
        RECT 96.630 119.210 96.800 119.380 ;
        RECT 98.300 120.650 98.470 120.820 ;
        RECT 98.300 120.290 98.470 120.460 ;
        RECT 98.300 119.930 98.470 120.100 ;
        RECT 98.300 119.570 98.470 119.740 ;
        RECT 98.300 119.210 98.470 119.380 ;
        RECT 100.220 120.650 100.390 120.820 ;
        RECT 100.220 120.290 100.390 120.460 ;
        RECT 100.220 119.930 100.390 120.100 ;
        RECT 100.220 119.570 100.390 119.740 ;
        RECT 100.220 119.210 100.390 119.380 ;
        RECT 102.440 120.550 102.610 120.720 ;
        RECT 102.440 120.190 102.610 120.360 ;
        RECT 102.440 119.830 102.610 120.000 ;
        RECT 102.440 119.470 102.610 119.640 ;
        RECT 102.440 119.110 102.610 119.280 ;
        RECT 96.080 118.750 96.250 118.920 ;
        RECT 97.285 118.790 97.455 118.960 ;
        RECT 97.645 118.790 97.815 118.960 ;
        RECT 100.875 118.790 101.045 118.960 ;
        RECT 101.235 118.790 101.405 118.960 ;
        RECT 96.080 118.390 96.250 118.560 ;
        RECT 102.440 118.750 102.610 118.920 ;
        RECT 96.080 118.030 96.250 118.200 ;
        RECT 96.080 117.670 96.250 117.840 ;
        RECT 86.030 117.230 86.200 117.400 ;
        RECT 86.030 116.870 86.200 117.040 ;
        RECT 82.740 116.245 82.910 116.415 ;
        RECT 86.030 116.510 86.200 116.680 ;
        RECT 84.895 116.230 85.065 116.400 ;
        RECT 82.740 115.885 82.910 116.055 ;
        RECT 86.030 116.150 86.200 116.320 ;
        RECT 82.740 115.525 82.910 115.695 ;
        RECT 82.740 115.165 82.910 115.335 ;
        RECT 82.740 114.805 82.910 114.975 ;
        RECT 82.740 114.445 82.910 114.615 ;
        RECT 84.310 115.845 84.480 116.015 ;
        RECT 84.310 115.485 84.480 115.655 ;
        RECT 84.310 115.125 84.480 115.295 ;
        RECT 86.030 115.790 86.200 115.960 ;
        RECT 86.030 115.430 86.200 115.600 ;
        RECT 84.895 114.950 85.065 115.120 ;
        RECT 86.030 115.070 86.200 115.240 ;
        RECT 84.310 114.765 84.480 114.935 ;
        RECT 84.310 114.405 84.480 114.575 ;
        RECT 81.020 113.990 81.190 114.160 ;
        RECT 82.155 114.070 82.325 114.240 ;
        RECT 84.310 114.045 84.480 114.215 ;
        RECT 86.030 114.710 86.200 114.880 ;
        RECT 86.030 114.350 86.200 114.520 ;
        RECT 86.030 113.990 86.200 114.160 ;
        RECT 81.020 113.630 81.190 113.800 ;
        RECT 84.895 113.670 85.065 113.840 ;
        RECT 86.030 113.630 86.200 113.800 ;
        RECT 96.080 117.310 96.250 117.480 ;
        RECT 96.080 116.950 96.250 117.120 ;
        RECT 96.630 118.370 96.800 118.540 ;
        RECT 96.630 118.010 96.800 118.180 ;
        RECT 96.630 117.650 96.800 117.820 ;
        RECT 96.630 117.290 96.800 117.460 ;
        RECT 96.630 116.930 96.800 117.100 ;
        RECT 98.300 118.370 98.470 118.540 ;
        RECT 98.300 118.010 98.470 118.180 ;
        RECT 98.300 117.650 98.470 117.820 ;
        RECT 98.300 117.290 98.470 117.460 ;
        RECT 98.300 116.930 98.470 117.100 ;
        RECT 100.220 118.370 100.390 118.540 ;
        RECT 100.220 118.010 100.390 118.180 ;
        RECT 100.220 117.650 100.390 117.820 ;
        RECT 100.220 117.290 100.390 117.460 ;
        RECT 100.220 116.930 100.390 117.100 ;
        RECT 102.440 118.390 102.610 118.560 ;
        RECT 102.440 118.030 102.610 118.200 ;
        RECT 102.440 117.670 102.610 117.840 ;
        RECT 102.440 117.310 102.610 117.480 ;
        RECT 102.440 116.950 102.610 117.120 ;
        RECT 96.080 116.590 96.250 116.760 ;
        RECT 97.285 116.510 97.455 116.680 ;
        RECT 97.645 116.510 97.815 116.680 ;
        RECT 100.875 116.510 101.045 116.680 ;
        RECT 101.235 116.510 101.405 116.680 ;
        RECT 102.440 116.590 102.610 116.760 ;
        RECT 96.080 116.230 96.250 116.400 ;
        RECT 96.080 115.870 96.250 116.040 ;
        RECT 96.080 115.510 96.250 115.680 ;
        RECT 96.080 115.150 96.250 115.320 ;
        RECT 96.080 114.790 96.250 114.960 ;
        RECT 96.630 116.090 96.800 116.260 ;
        RECT 96.630 115.730 96.800 115.900 ;
        RECT 96.630 115.370 96.800 115.540 ;
        RECT 96.630 115.010 96.800 115.180 ;
        RECT 96.630 114.650 96.800 114.820 ;
        RECT 98.300 116.090 98.470 116.260 ;
        RECT 98.300 115.730 98.470 115.900 ;
        RECT 98.300 115.370 98.470 115.540 ;
        RECT 98.300 115.010 98.470 115.180 ;
        RECT 98.300 114.650 98.470 114.820 ;
        RECT 100.220 116.090 100.390 116.260 ;
        RECT 100.220 115.730 100.390 115.900 ;
        RECT 100.220 115.370 100.390 115.540 ;
        RECT 100.220 115.010 100.390 115.180 ;
        RECT 100.220 114.650 100.390 114.820 ;
        RECT 102.440 116.230 102.610 116.400 ;
        RECT 102.440 115.870 102.610 116.040 ;
        RECT 102.440 115.510 102.610 115.680 ;
        RECT 102.440 115.150 102.610 115.320 ;
        RECT 102.440 114.790 102.610 114.960 ;
        RECT 96.080 114.430 96.250 114.600 ;
        RECT 102.440 114.430 102.610 114.600 ;
        RECT 96.080 114.070 96.250 114.240 ;
        RECT 97.285 114.230 97.455 114.400 ;
        RECT 97.645 114.230 97.815 114.400 ;
        RECT 100.875 114.230 101.045 114.400 ;
        RECT 101.235 114.230 101.405 114.400 ;
        RECT 102.440 114.070 102.610 114.240 ;
        RECT 96.080 113.710 96.250 113.880 ;
        RECT 98.300 113.810 98.470 113.980 ;
        RECT 81.320 113.040 81.490 113.210 ;
        RECT 81.680 113.040 81.850 113.210 ;
        RECT 82.040 113.040 82.210 113.210 ;
        RECT 82.400 113.040 82.570 113.210 ;
        RECT 82.760 113.040 82.930 113.210 ;
        RECT 83.120 113.040 83.290 113.210 ;
        RECT 83.480 113.040 83.650 113.210 ;
        RECT 83.840 113.040 84.010 113.210 ;
        RECT 84.200 113.040 84.370 113.210 ;
        RECT 84.560 113.040 84.730 113.210 ;
        RECT 84.920 113.040 85.090 113.210 ;
        RECT 85.280 113.040 85.450 113.210 ;
        RECT 85.640 113.040 85.810 113.210 ;
        RECT 88.845 113.340 89.015 113.510 ;
        RECT 89.205 113.340 89.375 113.510 ;
        RECT 89.565 113.340 89.735 113.510 ;
        RECT 89.925 113.340 90.095 113.510 ;
        RECT 90.285 113.340 90.455 113.510 ;
        RECT 90.645 113.340 90.815 113.510 ;
        RECT 92.115 113.340 92.285 113.510 ;
        RECT 92.475 113.340 92.645 113.510 ;
        RECT 92.835 113.340 93.005 113.510 ;
        RECT 93.195 113.340 93.365 113.510 ;
        RECT 93.555 113.340 93.725 113.510 ;
        RECT 93.915 113.340 94.085 113.510 ;
        RECT 94.275 113.340 94.445 113.510 ;
        RECT 94.635 113.340 94.805 113.510 ;
        RECT 63.685 112.630 63.855 112.800 ;
        RECT 64.550 112.670 64.720 112.840 ;
        RECT 64.910 112.670 65.080 112.840 ;
        RECT 69.280 112.670 69.450 112.840 ;
        RECT 63.685 112.270 63.855 112.440 ;
        RECT 70.075 112.630 70.245 112.800 ;
        RECT 63.685 111.910 63.855 112.080 ;
        RECT 63.685 111.550 63.855 111.720 ;
        RECT 63.685 111.190 63.855 111.360 ;
        RECT 63.685 110.830 63.855 111.000 ;
        RECT 65.565 112.250 65.735 112.420 ;
        RECT 65.565 111.890 65.735 112.060 ;
        RECT 65.565 111.530 65.735 111.700 ;
        RECT 65.565 111.170 65.735 111.340 ;
        RECT 65.565 110.810 65.735 110.980 ;
        RECT 68.695 112.250 68.865 112.420 ;
        RECT 68.695 111.890 68.865 112.060 ;
        RECT 68.695 111.530 68.865 111.700 ;
        RECT 68.695 111.170 68.865 111.340 ;
        RECT 68.695 110.810 68.865 110.980 ;
        RECT 70.075 112.270 70.245 112.440 ;
        RECT 70.075 111.910 70.245 112.080 ;
        RECT 70.075 111.550 70.245 111.720 ;
        RECT 70.075 111.190 70.245 111.360 ;
        RECT 70.075 110.830 70.245 111.000 ;
        RECT 63.685 110.470 63.855 110.640 ;
        RECT 64.550 110.390 64.720 110.560 ;
        RECT 64.910 110.390 65.080 110.560 ;
        RECT 69.280 110.390 69.450 110.560 ;
        RECT 70.075 110.470 70.245 110.640 ;
        RECT 63.685 110.110 63.855 110.280 ;
        RECT 63.685 109.750 63.855 109.920 ;
        RECT 63.685 109.390 63.855 109.560 ;
        RECT 63.685 109.030 63.855 109.200 ;
        RECT 63.685 108.670 63.855 108.840 ;
        RECT 65.565 109.970 65.735 110.140 ;
        RECT 65.565 109.610 65.735 109.780 ;
        RECT 65.565 109.250 65.735 109.420 ;
        RECT 65.565 108.890 65.735 109.060 ;
        RECT 65.565 108.530 65.735 108.700 ;
        RECT 68.695 109.970 68.865 110.140 ;
        RECT 68.695 109.610 68.865 109.780 ;
        RECT 68.695 109.250 68.865 109.420 ;
        RECT 68.695 108.890 68.865 109.060 ;
        RECT 68.695 108.530 68.865 108.700 ;
        RECT 70.075 110.110 70.245 110.280 ;
        RECT 70.075 109.750 70.245 109.920 ;
        RECT 70.075 109.390 70.245 109.560 ;
        RECT 70.075 109.030 70.245 109.200 ;
        RECT 70.075 108.670 70.245 108.840 ;
        RECT 63.685 108.310 63.855 108.480 ;
        RECT 70.075 108.310 70.245 108.480 ;
        RECT 63.685 107.950 63.855 108.120 ;
        RECT 64.550 108.110 64.720 108.280 ;
        RECT 64.910 108.110 65.080 108.280 ;
        RECT 69.280 108.110 69.450 108.280 ;
        RECT 70.075 107.950 70.245 108.120 ;
        RECT 63.685 107.590 63.855 107.760 ;
        RECT 63.685 107.230 63.855 107.400 ;
        RECT 63.685 106.870 63.855 107.040 ;
        RECT 63.685 106.510 63.855 106.680 ;
        RECT 63.685 106.150 63.855 106.320 ;
        RECT 65.565 107.690 65.735 107.860 ;
        RECT 65.565 107.330 65.735 107.500 ;
        RECT 65.565 106.970 65.735 107.140 ;
        RECT 65.565 106.610 65.735 106.780 ;
        RECT 65.565 106.250 65.735 106.420 ;
        RECT 68.695 107.690 68.865 107.860 ;
        RECT 68.695 107.330 68.865 107.500 ;
        RECT 68.695 106.970 68.865 107.140 ;
        RECT 68.695 106.610 68.865 106.780 ;
        RECT 68.695 106.250 68.865 106.420 ;
        RECT 70.075 107.590 70.245 107.760 ;
        RECT 70.075 107.230 70.245 107.400 ;
        RECT 70.075 106.870 70.245 107.040 ;
        RECT 70.075 106.510 70.245 106.680 ;
        RECT 70.075 106.150 70.245 106.320 ;
        RECT 63.685 105.790 63.855 105.960 ;
        RECT 64.550 105.830 64.720 106.000 ;
        RECT 64.910 105.830 65.080 106.000 ;
        RECT 69.280 105.830 69.450 106.000 ;
        RECT 63.685 105.430 63.855 105.600 ;
        RECT 70.075 105.790 70.245 105.960 ;
        RECT 63.685 105.070 63.855 105.240 ;
        RECT 63.685 104.710 63.855 104.880 ;
        RECT 63.685 104.350 63.855 104.520 ;
        RECT 63.685 103.990 63.855 104.160 ;
        RECT 65.565 105.410 65.735 105.580 ;
        RECT 65.565 105.050 65.735 105.220 ;
        RECT 65.565 104.690 65.735 104.860 ;
        RECT 65.565 104.330 65.735 104.500 ;
        RECT 65.565 103.970 65.735 104.140 ;
        RECT 68.695 105.410 68.865 105.580 ;
        RECT 68.695 105.050 68.865 105.220 ;
        RECT 68.695 104.690 68.865 104.860 ;
        RECT 68.695 104.330 68.865 104.500 ;
        RECT 68.695 103.970 68.865 104.140 ;
        RECT 70.075 105.430 70.245 105.600 ;
        RECT 70.075 105.070 70.245 105.240 ;
        RECT 70.075 104.710 70.245 104.880 ;
        RECT 70.075 104.350 70.245 104.520 ;
        RECT 70.075 103.990 70.245 104.160 ;
        RECT 63.685 103.630 63.855 103.800 ;
        RECT 64.550 103.550 64.720 103.720 ;
        RECT 64.910 103.550 65.080 103.720 ;
        RECT 69.280 103.550 69.450 103.720 ;
        RECT 70.075 103.630 70.245 103.800 ;
        RECT 63.685 103.270 63.855 103.440 ;
        RECT 63.685 102.910 63.855 103.080 ;
        RECT 63.685 102.550 63.855 102.720 ;
        RECT 63.685 102.190 63.855 102.360 ;
        RECT 63.685 101.830 63.855 102.000 ;
        RECT 65.565 103.130 65.735 103.300 ;
        RECT 65.565 102.770 65.735 102.940 ;
        RECT 65.565 102.410 65.735 102.580 ;
        RECT 65.565 102.050 65.735 102.220 ;
        RECT 65.565 101.690 65.735 101.860 ;
        RECT 68.695 103.130 68.865 103.300 ;
        RECT 68.695 102.770 68.865 102.940 ;
        RECT 68.695 102.410 68.865 102.580 ;
        RECT 68.695 102.050 68.865 102.220 ;
        RECT 68.695 101.690 68.865 101.860 ;
        RECT 70.075 103.270 70.245 103.440 ;
        RECT 70.075 102.910 70.245 103.080 ;
        RECT 70.075 102.550 70.245 102.720 ;
        RECT 70.075 102.190 70.245 102.360 ;
        RECT 70.075 101.830 70.245 102.000 ;
        RECT 63.685 101.470 63.855 101.640 ;
        RECT 70.075 101.470 70.245 101.640 ;
        RECT 63.685 101.110 63.855 101.280 ;
        RECT 64.550 101.270 64.720 101.440 ;
        RECT 64.910 101.270 65.080 101.440 ;
        RECT 69.280 101.270 69.450 101.440 ;
        RECT 70.075 101.110 70.245 101.280 ;
        RECT 63.685 100.750 63.855 100.920 ;
        RECT 63.685 100.390 63.855 100.560 ;
        RECT 63.685 100.030 63.855 100.200 ;
        RECT 63.685 99.670 63.855 99.840 ;
        RECT 63.685 99.310 63.855 99.480 ;
        RECT 65.565 100.850 65.735 101.020 ;
        RECT 65.565 100.490 65.735 100.660 ;
        RECT 65.565 100.130 65.735 100.300 ;
        RECT 65.565 99.770 65.735 99.940 ;
        RECT 65.565 99.410 65.735 99.580 ;
        RECT 68.695 100.850 68.865 101.020 ;
        RECT 68.695 100.490 68.865 100.660 ;
        RECT 68.695 100.130 68.865 100.300 ;
        RECT 68.695 99.770 68.865 99.940 ;
        RECT 68.695 99.410 68.865 99.580 ;
        RECT 70.075 100.750 70.245 100.920 ;
        RECT 70.075 100.390 70.245 100.560 ;
        RECT 70.075 100.030 70.245 100.200 ;
        RECT 70.075 99.670 70.245 99.840 ;
        RECT 70.075 99.310 70.245 99.480 ;
        RECT 63.685 98.950 63.855 99.120 ;
        RECT 64.550 98.990 64.720 99.160 ;
        RECT 64.910 98.990 65.080 99.160 ;
        RECT 69.280 98.990 69.450 99.160 ;
        RECT 63.685 98.590 63.855 98.760 ;
        RECT 70.075 98.950 70.245 99.120 ;
        RECT 63.685 98.230 63.855 98.400 ;
        RECT 63.685 97.870 63.855 98.040 ;
        RECT 63.685 97.510 63.855 97.680 ;
        RECT 63.685 97.150 63.855 97.320 ;
        RECT 65.565 98.570 65.735 98.740 ;
        RECT 65.565 98.210 65.735 98.380 ;
        RECT 65.565 97.850 65.735 98.020 ;
        RECT 65.565 97.490 65.735 97.660 ;
        RECT 65.565 97.130 65.735 97.300 ;
        RECT 68.695 98.570 68.865 98.740 ;
        RECT 68.695 98.210 68.865 98.380 ;
        RECT 68.695 97.850 68.865 98.020 ;
        RECT 68.695 97.490 68.865 97.660 ;
        RECT 68.695 97.130 68.865 97.300 ;
        RECT 70.075 98.590 70.245 98.760 ;
        RECT 70.075 98.230 70.245 98.400 ;
        RECT 70.075 97.870 70.245 98.040 ;
        RECT 70.075 97.510 70.245 97.680 ;
        RECT 70.075 97.150 70.245 97.320 ;
        RECT 63.685 96.790 63.855 96.960 ;
        RECT 64.550 96.710 64.720 96.880 ;
        RECT 64.910 96.710 65.080 96.880 ;
        RECT 69.280 96.710 69.450 96.880 ;
        RECT 70.075 96.790 70.245 96.960 ;
        RECT 63.685 96.430 63.855 96.600 ;
        RECT 63.685 96.070 63.855 96.240 ;
        RECT 63.685 95.710 63.855 95.880 ;
        RECT 63.685 95.350 63.855 95.520 ;
        RECT 63.685 94.990 63.855 95.160 ;
        RECT 65.565 96.290 65.735 96.460 ;
        RECT 65.565 95.930 65.735 96.100 ;
        RECT 65.565 95.570 65.735 95.740 ;
        RECT 65.565 95.210 65.735 95.380 ;
        RECT 65.565 94.850 65.735 95.020 ;
        RECT 68.695 96.290 68.865 96.460 ;
        RECT 68.695 95.930 68.865 96.100 ;
        RECT 68.695 95.570 68.865 95.740 ;
        RECT 68.695 95.210 68.865 95.380 ;
        RECT 68.695 94.850 68.865 95.020 ;
        RECT 70.075 96.430 70.245 96.600 ;
        RECT 70.075 96.070 70.245 96.240 ;
        RECT 70.075 95.710 70.245 95.880 ;
        RECT 70.075 95.350 70.245 95.520 ;
        RECT 70.075 94.990 70.245 95.160 ;
        RECT 63.685 94.630 63.855 94.800 ;
        RECT 70.075 94.630 70.245 94.800 ;
        RECT 63.685 94.270 63.855 94.440 ;
        RECT 64.550 94.430 64.720 94.600 ;
        RECT 64.910 94.430 65.080 94.600 ;
        RECT 69.280 94.430 69.450 94.600 ;
        RECT 70.075 94.270 70.245 94.440 ;
        RECT 63.685 93.910 63.855 94.080 ;
        RECT 63.685 93.550 63.855 93.720 ;
        RECT 63.685 93.190 63.855 93.360 ;
        RECT 63.685 92.830 63.855 93.000 ;
        RECT 63.685 92.470 63.855 92.640 ;
        RECT 65.565 94.010 65.735 94.180 ;
        RECT 65.565 93.650 65.735 93.820 ;
        RECT 65.565 93.290 65.735 93.460 ;
        RECT 65.565 92.930 65.735 93.100 ;
        RECT 65.565 92.570 65.735 92.740 ;
        RECT 68.695 94.010 68.865 94.180 ;
        RECT 68.695 93.650 68.865 93.820 ;
        RECT 68.695 93.290 68.865 93.460 ;
        RECT 68.695 92.930 68.865 93.100 ;
        RECT 68.695 92.570 68.865 92.740 ;
        RECT 70.075 93.910 70.245 94.080 ;
        RECT 70.075 93.550 70.245 93.720 ;
        RECT 70.075 93.190 70.245 93.360 ;
        RECT 70.075 92.830 70.245 93.000 ;
        RECT 70.075 92.470 70.245 92.640 ;
        RECT 63.685 92.110 63.855 92.280 ;
        RECT 64.550 92.150 64.720 92.320 ;
        RECT 64.910 92.150 65.080 92.320 ;
        RECT 69.280 92.150 69.450 92.320 ;
        RECT 63.685 91.750 63.855 91.920 ;
        RECT 70.075 92.110 70.245 92.280 ;
        RECT 63.685 91.390 63.855 91.560 ;
        RECT 63.685 91.030 63.855 91.200 ;
        RECT 63.685 90.670 63.855 90.840 ;
        RECT 63.685 90.310 63.855 90.480 ;
        RECT 65.565 91.730 65.735 91.900 ;
        RECT 65.565 91.370 65.735 91.540 ;
        RECT 65.565 91.010 65.735 91.180 ;
        RECT 65.565 90.650 65.735 90.820 ;
        RECT 65.565 90.290 65.735 90.460 ;
        RECT 68.695 91.730 68.865 91.900 ;
        RECT 68.695 91.370 68.865 91.540 ;
        RECT 68.695 91.010 68.865 91.180 ;
        RECT 68.695 90.650 68.865 90.820 ;
        RECT 68.695 90.290 68.865 90.460 ;
        RECT 70.075 91.750 70.245 91.920 ;
        RECT 70.075 91.390 70.245 91.560 ;
        RECT 70.075 91.030 70.245 91.200 ;
        RECT 70.075 90.670 70.245 90.840 ;
        RECT 70.075 90.310 70.245 90.480 ;
        RECT 63.685 89.950 63.855 90.120 ;
        RECT 64.550 89.870 64.720 90.040 ;
        RECT 64.910 89.870 65.080 90.040 ;
        RECT 69.280 89.870 69.450 90.040 ;
        RECT 70.075 89.950 70.245 90.120 ;
        RECT 63.685 89.590 63.855 89.760 ;
        RECT 70.075 89.590 70.245 89.760 ;
        RECT 63.985 89.200 64.155 89.370 ;
        RECT 64.345 89.200 64.515 89.370 ;
        RECT 64.705 89.200 64.875 89.370 ;
        RECT 65.065 89.200 65.235 89.370 ;
        RECT 65.425 89.200 65.595 89.370 ;
        RECT 65.785 89.200 65.955 89.370 ;
        RECT 66.145 89.200 66.315 89.370 ;
        RECT 66.505 89.200 66.675 89.370 ;
        RECT 67.975 89.200 68.145 89.370 ;
        RECT 68.335 89.200 68.505 89.370 ;
        RECT 68.695 89.200 68.865 89.370 ;
        RECT 69.055 89.200 69.225 89.370 ;
        RECT 69.415 89.200 69.585 89.370 ;
        RECT 69.775 89.200 69.945 89.370 ;
        RECT 88.545 112.990 88.715 113.160 ;
        RECT 94.935 112.990 95.105 113.160 ;
        RECT 88.545 112.630 88.715 112.800 ;
        RECT 89.340 112.670 89.510 112.840 ;
        RECT 93.710 112.670 93.880 112.840 ;
        RECT 94.070 112.670 94.240 112.840 ;
        RECT 88.545 112.270 88.715 112.440 ;
        RECT 94.935 112.630 95.105 112.800 ;
        RECT 88.545 111.910 88.715 112.080 ;
        RECT 88.545 111.550 88.715 111.720 ;
        RECT 88.545 111.190 88.715 111.360 ;
        RECT 88.545 110.830 88.715 111.000 ;
        RECT 89.925 112.250 90.095 112.420 ;
        RECT 89.925 111.890 90.095 112.060 ;
        RECT 89.925 111.530 90.095 111.700 ;
        RECT 89.925 111.170 90.095 111.340 ;
        RECT 89.925 110.810 90.095 110.980 ;
        RECT 93.055 112.250 93.225 112.420 ;
        RECT 93.055 111.890 93.225 112.060 ;
        RECT 93.055 111.530 93.225 111.700 ;
        RECT 93.055 111.170 93.225 111.340 ;
        RECT 93.055 110.810 93.225 110.980 ;
        RECT 94.935 112.270 95.105 112.440 ;
        RECT 94.935 111.910 95.105 112.080 ;
        RECT 96.080 113.350 96.250 113.520 ;
        RECT 97.285 113.450 97.455 113.620 ;
        RECT 97.645 113.450 97.815 113.620 ;
        RECT 98.300 113.450 98.470 113.620 ;
        RECT 96.080 112.990 96.250 113.160 ;
        RECT 98.300 113.090 98.470 113.260 ;
        RECT 102.440 113.710 102.610 113.880 ;
        RECT 102.440 113.350 102.610 113.520 ;
        RECT 102.440 112.990 102.610 113.160 ;
        RECT 96.080 112.630 96.250 112.800 ;
        RECT 97.285 112.670 97.455 112.840 ;
        RECT 97.645 112.670 97.815 112.840 ;
        RECT 102.440 112.630 102.610 112.800 ;
        RECT 96.380 112.000 96.550 112.170 ;
        RECT 96.740 112.000 96.910 112.170 ;
        RECT 97.100 112.000 97.270 112.170 ;
        RECT 97.460 112.000 97.630 112.170 ;
        RECT 97.820 112.000 97.990 112.170 ;
        RECT 98.180 112.000 98.350 112.170 ;
        RECT 98.540 112.000 98.710 112.170 ;
        RECT 98.900 112.000 99.070 112.170 ;
        RECT 99.260 112.000 99.430 112.170 ;
        RECT 99.620 112.000 99.790 112.170 ;
        RECT 99.980 112.000 100.150 112.170 ;
        RECT 100.340 112.000 100.510 112.170 ;
        RECT 100.700 112.000 100.870 112.170 ;
        RECT 101.060 112.000 101.230 112.170 ;
        RECT 101.420 112.000 101.590 112.170 ;
        RECT 101.780 112.000 101.950 112.170 ;
        RECT 102.140 112.000 102.310 112.170 ;
        RECT 108.635 151.370 108.805 151.540 ;
        RECT 108.635 151.010 108.805 151.180 ;
        RECT 110.555 152.260 110.725 152.430 ;
        RECT 110.555 151.900 110.725 152.070 ;
        RECT 110.555 151.540 110.725 151.710 ;
        RECT 110.555 151.180 110.725 151.350 ;
        RECT 110.555 150.820 110.725 150.990 ;
        RECT 111.925 152.260 112.095 152.430 ;
        RECT 111.925 151.900 112.095 152.070 ;
        RECT 111.925 151.540 112.095 151.710 ;
        RECT 111.925 151.180 112.095 151.350 ;
        RECT 111.925 150.820 112.095 150.990 ;
        RECT 113.845 152.070 114.015 152.240 ;
        RECT 113.845 151.710 114.015 151.880 ;
        RECT 113.845 151.350 114.015 151.520 ;
        RECT 113.845 150.990 114.015 151.160 ;
        RECT 108.635 150.650 108.805 150.820 ;
        RECT 113.845 150.630 114.015 150.800 ;
        RECT 108.635 150.290 108.805 150.460 ;
        RECT 109.690 150.400 109.860 150.570 ;
        RECT 110.050 150.400 110.220 150.570 ;
        RECT 111.060 150.400 111.230 150.570 ;
        RECT 111.420 150.400 111.590 150.570 ;
        RECT 112.430 150.400 112.600 150.570 ;
        RECT 112.790 150.400 112.960 150.570 ;
        RECT 113.845 150.270 114.015 150.440 ;
        RECT 108.635 149.930 108.805 150.100 ;
        RECT 108.635 149.570 108.805 149.740 ;
        RECT 108.635 149.210 108.805 149.380 ;
        RECT 108.635 148.850 108.805 149.020 ;
        RECT 108.635 148.490 108.805 148.660 ;
        RECT 110.555 149.980 110.725 150.150 ;
        RECT 110.555 149.620 110.725 149.790 ;
        RECT 110.555 149.260 110.725 149.430 ;
        RECT 110.555 148.900 110.725 149.070 ;
        RECT 110.555 148.540 110.725 148.710 ;
        RECT 111.925 149.980 112.095 150.150 ;
        RECT 111.925 149.620 112.095 149.790 ;
        RECT 111.925 149.260 112.095 149.430 ;
        RECT 111.925 148.900 112.095 149.070 ;
        RECT 111.925 148.540 112.095 148.710 ;
        RECT 113.845 149.910 114.015 150.080 ;
        RECT 113.845 149.550 114.015 149.720 ;
        RECT 113.845 149.190 114.015 149.360 ;
        RECT 113.845 148.830 114.015 149.000 ;
        RECT 108.635 148.130 108.805 148.300 ;
        RECT 113.845 148.470 114.015 148.640 ;
        RECT 109.690 148.120 109.860 148.290 ;
        RECT 110.050 148.120 110.220 148.290 ;
        RECT 111.060 148.120 111.230 148.290 ;
        RECT 111.420 148.120 111.590 148.290 ;
        RECT 112.430 148.120 112.600 148.290 ;
        RECT 112.790 148.120 112.960 148.290 ;
        RECT 108.635 147.770 108.805 147.940 ;
        RECT 113.845 148.110 114.015 148.280 ;
        RECT 108.635 147.410 108.805 147.580 ;
        RECT 108.635 147.050 108.805 147.220 ;
        RECT 108.635 146.690 108.805 146.860 ;
        RECT 108.635 146.330 108.805 146.500 ;
        RECT 110.555 147.700 110.725 147.870 ;
        RECT 110.555 147.340 110.725 147.510 ;
        RECT 110.555 146.980 110.725 147.150 ;
        RECT 110.555 146.620 110.725 146.790 ;
        RECT 110.555 146.260 110.725 146.430 ;
        RECT 111.925 147.700 112.095 147.870 ;
        RECT 111.925 147.340 112.095 147.510 ;
        RECT 111.925 146.980 112.095 147.150 ;
        RECT 111.925 146.620 112.095 146.790 ;
        RECT 111.925 146.260 112.095 146.430 ;
        RECT 113.845 147.750 114.015 147.920 ;
        RECT 113.845 147.390 114.015 147.560 ;
        RECT 113.845 147.030 114.015 147.200 ;
        RECT 113.845 146.670 114.015 146.840 ;
        RECT 113.845 146.310 114.015 146.480 ;
        RECT 108.635 145.970 108.805 146.140 ;
        RECT 109.690 145.840 109.860 146.010 ;
        RECT 110.050 145.840 110.220 146.010 ;
        RECT 111.060 145.840 111.230 146.010 ;
        RECT 111.420 145.840 111.590 146.010 ;
        RECT 112.430 145.840 112.600 146.010 ;
        RECT 112.790 145.840 112.960 146.010 ;
        RECT 113.845 145.950 114.015 146.120 ;
        RECT 108.635 145.610 108.805 145.780 ;
        RECT 113.845 145.590 114.015 145.760 ;
        RECT 108.635 145.250 108.805 145.420 ;
        RECT 108.635 144.890 108.805 145.060 ;
        RECT 108.635 144.530 108.805 144.700 ;
        RECT 108.635 144.170 108.805 144.340 ;
        RECT 110.555 145.420 110.725 145.590 ;
        RECT 110.555 145.060 110.725 145.230 ;
        RECT 110.555 144.700 110.725 144.870 ;
        RECT 110.555 144.340 110.725 144.510 ;
        RECT 110.555 143.980 110.725 144.150 ;
        RECT 111.925 145.420 112.095 145.590 ;
        RECT 111.925 145.060 112.095 145.230 ;
        RECT 111.925 144.700 112.095 144.870 ;
        RECT 111.925 144.340 112.095 144.510 ;
        RECT 111.925 143.980 112.095 144.150 ;
        RECT 113.845 145.230 114.015 145.400 ;
        RECT 113.845 144.870 114.015 145.040 ;
        RECT 113.845 144.510 114.015 144.680 ;
        RECT 113.845 144.150 114.015 144.320 ;
        RECT 108.635 143.810 108.805 143.980 ;
        RECT 113.845 143.790 114.015 143.960 ;
        RECT 108.635 143.450 108.805 143.620 ;
        RECT 109.690 143.560 109.860 143.730 ;
        RECT 110.050 143.560 110.220 143.730 ;
        RECT 111.060 143.560 111.230 143.730 ;
        RECT 111.420 143.560 111.590 143.730 ;
        RECT 112.430 143.560 112.600 143.730 ;
        RECT 112.790 143.560 112.960 143.730 ;
        RECT 113.845 143.430 114.015 143.600 ;
        RECT 108.635 143.090 108.805 143.260 ;
        RECT 108.635 142.730 108.805 142.900 ;
        RECT 108.635 142.370 108.805 142.540 ;
        RECT 108.635 142.010 108.805 142.180 ;
        RECT 108.635 141.650 108.805 141.820 ;
        RECT 110.555 143.140 110.725 143.310 ;
        RECT 110.555 142.780 110.725 142.950 ;
        RECT 110.555 142.420 110.725 142.590 ;
        RECT 110.555 142.060 110.725 142.230 ;
        RECT 110.555 141.700 110.725 141.870 ;
        RECT 111.925 143.140 112.095 143.310 ;
        RECT 111.925 142.780 112.095 142.950 ;
        RECT 111.925 142.420 112.095 142.590 ;
        RECT 111.925 142.060 112.095 142.230 ;
        RECT 111.925 141.700 112.095 141.870 ;
        RECT 113.845 143.070 114.015 143.240 ;
        RECT 113.845 142.710 114.015 142.880 ;
        RECT 113.845 142.350 114.015 142.520 ;
        RECT 113.845 141.990 114.015 142.160 ;
        RECT 108.635 141.290 108.805 141.460 ;
        RECT 113.845 141.630 114.015 141.800 ;
        RECT 109.690 141.280 109.860 141.450 ;
        RECT 110.050 141.280 110.220 141.450 ;
        RECT 111.060 141.280 111.230 141.450 ;
        RECT 111.420 141.280 111.590 141.450 ;
        RECT 112.430 141.280 112.600 141.450 ;
        RECT 112.790 141.280 112.960 141.450 ;
        RECT 108.635 140.930 108.805 141.100 ;
        RECT 113.845 141.270 114.015 141.440 ;
        RECT 108.635 140.570 108.805 140.740 ;
        RECT 108.635 140.210 108.805 140.380 ;
        RECT 108.635 139.850 108.805 140.020 ;
        RECT 108.635 139.490 108.805 139.660 ;
        RECT 110.555 140.860 110.725 141.030 ;
        RECT 110.555 140.500 110.725 140.670 ;
        RECT 110.555 140.140 110.725 140.310 ;
        RECT 110.555 139.780 110.725 139.950 ;
        RECT 110.555 139.420 110.725 139.590 ;
        RECT 111.925 140.860 112.095 141.030 ;
        RECT 111.925 140.500 112.095 140.670 ;
        RECT 111.925 140.140 112.095 140.310 ;
        RECT 111.925 139.780 112.095 139.950 ;
        RECT 111.925 139.420 112.095 139.590 ;
        RECT 113.845 140.910 114.015 141.080 ;
        RECT 113.845 140.550 114.015 140.720 ;
        RECT 113.845 140.190 114.015 140.360 ;
        RECT 113.845 139.830 114.015 140.000 ;
        RECT 113.845 139.470 114.015 139.640 ;
        RECT 108.635 139.130 108.805 139.300 ;
        RECT 109.690 139.000 109.860 139.170 ;
        RECT 110.050 139.000 110.220 139.170 ;
        RECT 111.060 139.000 111.230 139.170 ;
        RECT 111.420 139.000 111.590 139.170 ;
        RECT 112.430 139.000 112.600 139.170 ;
        RECT 112.790 139.000 112.960 139.170 ;
        RECT 113.845 139.110 114.015 139.280 ;
        RECT 108.635 138.770 108.805 138.940 ;
        RECT 113.845 138.750 114.015 138.920 ;
        RECT 108.635 138.410 108.805 138.580 ;
        RECT 108.635 138.050 108.805 138.220 ;
        RECT 108.635 137.690 108.805 137.860 ;
        RECT 108.635 137.330 108.805 137.500 ;
        RECT 110.555 138.580 110.725 138.750 ;
        RECT 110.555 138.220 110.725 138.390 ;
        RECT 110.555 137.860 110.725 138.030 ;
        RECT 110.555 137.500 110.725 137.670 ;
        RECT 110.555 137.140 110.725 137.310 ;
        RECT 111.925 138.580 112.095 138.750 ;
        RECT 111.925 138.220 112.095 138.390 ;
        RECT 111.925 137.860 112.095 138.030 ;
        RECT 111.925 137.500 112.095 137.670 ;
        RECT 111.925 137.140 112.095 137.310 ;
        RECT 113.845 138.390 114.015 138.560 ;
        RECT 113.845 138.030 114.015 138.200 ;
        RECT 113.845 137.670 114.015 137.840 ;
        RECT 113.845 137.310 114.015 137.480 ;
        RECT 108.635 136.970 108.805 137.140 ;
        RECT 113.845 136.950 114.015 137.120 ;
        RECT 108.635 136.610 108.805 136.780 ;
        RECT 109.690 136.720 109.860 136.890 ;
        RECT 110.050 136.720 110.220 136.890 ;
        RECT 111.060 136.720 111.230 136.890 ;
        RECT 111.420 136.720 111.590 136.890 ;
        RECT 112.430 136.720 112.600 136.890 ;
        RECT 112.790 136.720 112.960 136.890 ;
        RECT 113.845 136.590 114.015 136.760 ;
        RECT 108.635 136.250 108.805 136.420 ;
        RECT 108.635 135.890 108.805 136.060 ;
        RECT 108.635 135.530 108.805 135.700 ;
        RECT 108.635 135.170 108.805 135.340 ;
        RECT 108.635 134.810 108.805 134.980 ;
        RECT 110.555 136.300 110.725 136.470 ;
        RECT 110.555 135.940 110.725 136.110 ;
        RECT 110.555 135.580 110.725 135.750 ;
        RECT 110.555 135.220 110.725 135.390 ;
        RECT 110.555 134.860 110.725 135.030 ;
        RECT 111.925 136.300 112.095 136.470 ;
        RECT 111.925 135.940 112.095 136.110 ;
        RECT 111.925 135.580 112.095 135.750 ;
        RECT 111.925 135.220 112.095 135.390 ;
        RECT 111.925 134.860 112.095 135.030 ;
        RECT 113.845 136.230 114.015 136.400 ;
        RECT 113.845 135.870 114.015 136.040 ;
        RECT 113.845 135.510 114.015 135.680 ;
        RECT 113.845 135.150 114.015 135.320 ;
        RECT 108.635 134.450 108.805 134.620 ;
        RECT 113.845 134.790 114.015 134.960 ;
        RECT 109.690 134.440 109.860 134.610 ;
        RECT 110.050 134.440 110.220 134.610 ;
        RECT 111.060 134.440 111.230 134.610 ;
        RECT 111.420 134.440 111.590 134.610 ;
        RECT 112.430 134.440 112.600 134.610 ;
        RECT 112.790 134.440 112.960 134.610 ;
        RECT 108.635 134.090 108.805 134.260 ;
        RECT 113.845 134.430 114.015 134.600 ;
        RECT 108.635 133.730 108.805 133.900 ;
        RECT 108.635 133.370 108.805 133.540 ;
        RECT 108.635 133.010 108.805 133.180 ;
        RECT 108.635 132.650 108.805 132.820 ;
        RECT 110.555 134.020 110.725 134.190 ;
        RECT 110.555 133.660 110.725 133.830 ;
        RECT 110.555 133.300 110.725 133.470 ;
        RECT 110.555 132.940 110.725 133.110 ;
        RECT 110.555 132.580 110.725 132.750 ;
        RECT 111.925 134.020 112.095 134.190 ;
        RECT 111.925 133.660 112.095 133.830 ;
        RECT 111.925 133.300 112.095 133.470 ;
        RECT 111.925 132.940 112.095 133.110 ;
        RECT 111.925 132.580 112.095 132.750 ;
        RECT 113.845 134.070 114.015 134.240 ;
        RECT 113.845 133.710 114.015 133.880 ;
        RECT 113.845 133.350 114.015 133.520 ;
        RECT 113.845 132.990 114.015 133.160 ;
        RECT 113.845 132.630 114.015 132.800 ;
        RECT 108.635 132.290 108.805 132.460 ;
        RECT 109.690 132.160 109.860 132.330 ;
        RECT 110.050 132.160 110.220 132.330 ;
        RECT 111.060 132.160 111.230 132.330 ;
        RECT 111.420 132.160 111.590 132.330 ;
        RECT 112.430 132.160 112.600 132.330 ;
        RECT 112.790 132.160 112.960 132.330 ;
        RECT 113.845 132.270 114.015 132.440 ;
        RECT 108.635 131.930 108.805 132.100 ;
        RECT 113.845 131.910 114.015 132.080 ;
        RECT 108.635 131.570 108.805 131.740 ;
        RECT 108.635 131.210 108.805 131.380 ;
        RECT 108.635 130.850 108.805 131.020 ;
        RECT 108.635 130.490 108.805 130.660 ;
        RECT 110.555 131.740 110.725 131.910 ;
        RECT 110.555 131.380 110.725 131.550 ;
        RECT 110.555 131.020 110.725 131.190 ;
        RECT 110.555 130.660 110.725 130.830 ;
        RECT 110.555 130.300 110.725 130.470 ;
        RECT 111.925 131.740 112.095 131.910 ;
        RECT 111.925 131.380 112.095 131.550 ;
        RECT 111.925 131.020 112.095 131.190 ;
        RECT 111.925 130.660 112.095 130.830 ;
        RECT 111.925 130.300 112.095 130.470 ;
        RECT 113.845 131.550 114.015 131.720 ;
        RECT 113.845 131.190 114.015 131.360 ;
        RECT 113.845 130.830 114.015 131.000 ;
        RECT 113.845 130.470 114.015 130.640 ;
        RECT 108.635 130.130 108.805 130.300 ;
        RECT 113.845 130.110 114.015 130.280 ;
        RECT 108.635 129.770 108.805 129.940 ;
        RECT 109.690 129.880 109.860 130.050 ;
        RECT 110.050 129.880 110.220 130.050 ;
        RECT 111.060 129.880 111.230 130.050 ;
        RECT 111.420 129.880 111.590 130.050 ;
        RECT 112.430 129.880 112.600 130.050 ;
        RECT 112.790 129.880 112.960 130.050 ;
        RECT 113.845 129.750 114.015 129.920 ;
        RECT 108.635 129.410 108.805 129.580 ;
        RECT 108.635 129.050 108.805 129.220 ;
        RECT 108.635 128.690 108.805 128.860 ;
        RECT 108.635 128.330 108.805 128.500 ;
        RECT 108.635 127.970 108.805 128.140 ;
        RECT 110.555 129.460 110.725 129.630 ;
        RECT 110.555 129.100 110.725 129.270 ;
        RECT 110.555 128.740 110.725 128.910 ;
        RECT 110.555 128.380 110.725 128.550 ;
        RECT 110.555 128.020 110.725 128.190 ;
        RECT 111.925 129.460 112.095 129.630 ;
        RECT 111.925 129.100 112.095 129.270 ;
        RECT 111.925 128.740 112.095 128.910 ;
        RECT 111.925 128.380 112.095 128.550 ;
        RECT 111.925 128.020 112.095 128.190 ;
        RECT 113.845 129.390 114.015 129.560 ;
        RECT 113.845 129.030 114.015 129.200 ;
        RECT 113.845 128.670 114.015 128.840 ;
        RECT 113.845 128.310 114.015 128.480 ;
        RECT 108.635 127.610 108.805 127.780 ;
        RECT 113.845 127.950 114.015 128.120 ;
        RECT 109.690 127.600 109.860 127.770 ;
        RECT 110.050 127.600 110.220 127.770 ;
        RECT 111.060 127.600 111.230 127.770 ;
        RECT 111.420 127.600 111.590 127.770 ;
        RECT 112.430 127.600 112.600 127.770 ;
        RECT 112.790 127.600 112.960 127.770 ;
        RECT 108.635 127.250 108.805 127.420 ;
        RECT 113.845 127.590 114.015 127.760 ;
        RECT 108.635 126.890 108.805 127.060 ;
        RECT 108.635 126.530 108.805 126.700 ;
        RECT 108.635 126.170 108.805 126.340 ;
        RECT 108.635 125.810 108.805 125.980 ;
        RECT 110.555 127.180 110.725 127.350 ;
        RECT 110.555 126.820 110.725 126.990 ;
        RECT 110.555 126.460 110.725 126.630 ;
        RECT 110.555 126.100 110.725 126.270 ;
        RECT 110.555 125.740 110.725 125.910 ;
        RECT 111.925 127.180 112.095 127.350 ;
        RECT 111.925 126.820 112.095 126.990 ;
        RECT 111.925 126.460 112.095 126.630 ;
        RECT 111.925 126.100 112.095 126.270 ;
        RECT 111.925 125.740 112.095 125.910 ;
        RECT 113.845 127.230 114.015 127.400 ;
        RECT 113.845 126.870 114.015 127.040 ;
        RECT 113.845 126.510 114.015 126.680 ;
        RECT 113.845 126.150 114.015 126.320 ;
        RECT 113.845 125.790 114.015 125.960 ;
        RECT 108.635 125.450 108.805 125.620 ;
        RECT 109.690 125.320 109.860 125.490 ;
        RECT 110.050 125.320 110.220 125.490 ;
        RECT 111.060 125.320 111.230 125.490 ;
        RECT 111.420 125.320 111.590 125.490 ;
        RECT 112.430 125.320 112.600 125.490 ;
        RECT 112.790 125.320 112.960 125.490 ;
        RECT 113.845 125.430 114.015 125.600 ;
        RECT 108.635 125.090 108.805 125.260 ;
        RECT 113.845 125.070 114.015 125.240 ;
        RECT 108.635 124.730 108.805 124.900 ;
        RECT 108.635 124.370 108.805 124.540 ;
        RECT 108.635 124.010 108.805 124.180 ;
        RECT 108.635 123.650 108.805 123.820 ;
        RECT 110.555 124.900 110.725 125.070 ;
        RECT 110.555 124.540 110.725 124.710 ;
        RECT 110.555 124.180 110.725 124.350 ;
        RECT 110.555 123.820 110.725 123.990 ;
        RECT 110.555 123.460 110.725 123.630 ;
        RECT 111.925 124.900 112.095 125.070 ;
        RECT 111.925 124.540 112.095 124.710 ;
        RECT 111.925 124.180 112.095 124.350 ;
        RECT 111.925 123.820 112.095 123.990 ;
        RECT 111.925 123.460 112.095 123.630 ;
        RECT 113.845 124.710 114.015 124.880 ;
        RECT 113.845 124.350 114.015 124.520 ;
        RECT 113.845 123.990 114.015 124.160 ;
        RECT 113.845 123.630 114.015 123.800 ;
        RECT 108.635 123.290 108.805 123.460 ;
        RECT 113.845 123.270 114.015 123.440 ;
        RECT 108.635 122.930 108.805 123.100 ;
        RECT 109.690 123.040 109.860 123.210 ;
        RECT 110.050 123.040 110.220 123.210 ;
        RECT 111.060 123.040 111.230 123.210 ;
        RECT 111.420 123.040 111.590 123.210 ;
        RECT 112.430 123.040 112.600 123.210 ;
        RECT 112.790 123.040 112.960 123.210 ;
        RECT 113.845 122.910 114.015 123.080 ;
        RECT 108.635 122.570 108.805 122.740 ;
        RECT 108.635 122.210 108.805 122.380 ;
        RECT 108.635 121.850 108.805 122.020 ;
        RECT 108.635 121.490 108.805 121.660 ;
        RECT 108.635 121.130 108.805 121.300 ;
        RECT 110.555 122.620 110.725 122.790 ;
        RECT 110.555 122.260 110.725 122.430 ;
        RECT 110.555 121.900 110.725 122.070 ;
        RECT 110.555 121.540 110.725 121.710 ;
        RECT 110.555 121.180 110.725 121.350 ;
        RECT 111.925 122.620 112.095 122.790 ;
        RECT 111.925 122.260 112.095 122.430 ;
        RECT 111.925 121.900 112.095 122.070 ;
        RECT 111.925 121.540 112.095 121.710 ;
        RECT 111.925 121.180 112.095 121.350 ;
        RECT 113.845 122.550 114.015 122.720 ;
        RECT 113.845 122.190 114.015 122.360 ;
        RECT 113.845 121.830 114.015 122.000 ;
        RECT 113.845 121.470 114.015 121.640 ;
        RECT 108.635 120.770 108.805 120.940 ;
        RECT 113.845 121.110 114.015 121.280 ;
        RECT 109.690 120.760 109.860 120.930 ;
        RECT 110.050 120.760 110.220 120.930 ;
        RECT 111.060 120.760 111.230 120.930 ;
        RECT 111.420 120.760 111.590 120.930 ;
        RECT 112.430 120.760 112.600 120.930 ;
        RECT 112.790 120.760 112.960 120.930 ;
        RECT 108.635 120.410 108.805 120.580 ;
        RECT 113.845 120.750 114.015 120.920 ;
        RECT 108.635 120.050 108.805 120.220 ;
        RECT 108.635 119.690 108.805 119.860 ;
        RECT 108.635 119.330 108.805 119.500 ;
        RECT 108.635 118.970 108.805 119.140 ;
        RECT 110.555 120.340 110.725 120.510 ;
        RECT 110.555 119.980 110.725 120.150 ;
        RECT 110.555 119.620 110.725 119.790 ;
        RECT 110.555 119.260 110.725 119.430 ;
        RECT 110.555 118.900 110.725 119.070 ;
        RECT 111.925 120.340 112.095 120.510 ;
        RECT 111.925 119.980 112.095 120.150 ;
        RECT 111.925 119.620 112.095 119.790 ;
        RECT 111.925 119.260 112.095 119.430 ;
        RECT 111.925 118.900 112.095 119.070 ;
        RECT 113.845 120.390 114.015 120.560 ;
        RECT 113.845 120.030 114.015 120.200 ;
        RECT 113.845 119.670 114.015 119.840 ;
        RECT 113.845 119.310 114.015 119.480 ;
        RECT 113.845 118.950 114.015 119.120 ;
        RECT 108.635 118.610 108.805 118.780 ;
        RECT 109.690 118.480 109.860 118.650 ;
        RECT 110.050 118.480 110.220 118.650 ;
        RECT 111.060 118.480 111.230 118.650 ;
        RECT 111.420 118.480 111.590 118.650 ;
        RECT 112.430 118.480 112.600 118.650 ;
        RECT 112.790 118.480 112.960 118.650 ;
        RECT 113.845 118.590 114.015 118.760 ;
        RECT 108.635 118.250 108.805 118.420 ;
        RECT 113.845 118.230 114.015 118.400 ;
        RECT 121.840 164.650 122.010 164.820 ;
        RECT 122.380 164.710 122.550 164.880 ;
        RECT 122.740 164.710 122.910 164.880 ;
        RECT 123.100 164.710 123.270 164.880 ;
        RECT 123.460 164.710 123.630 164.880 ;
        RECT 123.820 164.710 123.990 164.880 ;
        RECT 124.180 164.710 124.350 164.880 ;
        RECT 124.540 164.710 124.710 164.880 ;
        RECT 124.900 164.710 125.070 164.880 ;
        RECT 125.260 164.710 125.430 164.880 ;
        RECT 125.620 164.710 125.790 164.880 ;
        RECT 121.840 164.290 122.010 164.460 ;
        RECT 125.680 164.350 125.850 164.520 ;
        RECT 121.840 163.930 122.010 164.100 ;
        RECT 122.895 164.080 123.065 164.250 ;
        RECT 123.255 164.080 123.425 164.250 ;
        RECT 124.265 164.080 124.435 164.250 ;
        RECT 124.625 164.080 124.795 164.250 ;
        RECT 125.680 163.990 125.850 164.160 ;
        RECT 121.840 163.570 122.010 163.740 ;
        RECT 121.840 163.210 122.010 163.380 ;
        RECT 121.840 162.850 122.010 163.020 ;
        RECT 121.840 162.490 122.010 162.660 ;
        RECT 121.840 162.130 122.010 162.300 ;
        RECT 122.390 163.660 122.560 163.830 ;
        RECT 122.390 163.300 122.560 163.470 ;
        RECT 122.390 162.940 122.560 163.110 ;
        RECT 122.390 162.580 122.560 162.750 ;
        RECT 122.390 162.220 122.560 162.390 ;
        RECT 125.130 163.660 125.300 163.830 ;
        RECT 125.130 163.300 125.300 163.470 ;
        RECT 125.130 162.940 125.300 163.110 ;
        RECT 125.130 162.580 125.300 162.750 ;
        RECT 125.130 162.220 125.300 162.390 ;
        RECT 125.680 163.630 125.850 163.800 ;
        RECT 125.680 163.270 125.850 163.440 ;
        RECT 125.680 162.910 125.850 163.080 ;
        RECT 125.680 162.550 125.850 162.720 ;
        RECT 125.680 162.190 125.850 162.360 ;
        RECT 121.840 161.770 122.010 161.940 ;
        RECT 122.895 161.800 123.065 161.970 ;
        RECT 123.255 161.800 123.425 161.970 ;
        RECT 124.265 161.800 124.435 161.970 ;
        RECT 124.625 161.800 124.795 161.970 ;
        RECT 125.680 161.830 125.850 162.000 ;
        RECT 121.840 161.410 122.010 161.580 ;
        RECT 121.840 161.050 122.010 161.220 ;
        RECT 121.840 160.690 122.010 160.860 ;
        RECT 121.840 160.330 122.010 160.500 ;
        RECT 121.840 159.970 122.010 160.140 ;
        RECT 122.390 161.380 122.560 161.550 ;
        RECT 122.390 161.020 122.560 161.190 ;
        RECT 122.390 160.660 122.560 160.830 ;
        RECT 122.390 160.300 122.560 160.470 ;
        RECT 122.390 159.940 122.560 160.110 ;
        RECT 125.130 161.380 125.300 161.550 ;
        RECT 125.130 161.020 125.300 161.190 ;
        RECT 125.130 160.660 125.300 160.830 ;
        RECT 125.130 160.300 125.300 160.470 ;
        RECT 125.130 159.940 125.300 160.110 ;
        RECT 125.680 161.470 125.850 161.640 ;
        RECT 125.680 161.110 125.850 161.280 ;
        RECT 125.680 160.750 125.850 160.920 ;
        RECT 125.680 160.390 125.850 160.560 ;
        RECT 125.680 160.030 125.850 160.200 ;
        RECT 121.840 159.610 122.010 159.780 ;
        RECT 122.895 159.520 123.065 159.690 ;
        RECT 123.255 159.520 123.425 159.690 ;
        RECT 124.265 159.520 124.435 159.690 ;
        RECT 124.625 159.520 124.795 159.690 ;
        RECT 125.680 159.670 125.850 159.840 ;
        RECT 121.840 159.250 122.010 159.420 ;
        RECT 125.680 159.310 125.850 159.480 ;
        RECT 121.840 158.890 122.010 159.060 ;
        RECT 121.840 158.530 122.010 158.700 ;
        RECT 121.840 158.170 122.010 158.340 ;
        RECT 121.840 157.810 122.010 157.980 ;
        RECT 122.390 159.100 122.560 159.270 ;
        RECT 122.390 158.740 122.560 158.910 ;
        RECT 122.390 158.380 122.560 158.550 ;
        RECT 122.390 158.020 122.560 158.190 ;
        RECT 122.390 157.660 122.560 157.830 ;
        RECT 123.760 159.100 123.930 159.270 ;
        RECT 123.760 158.740 123.930 158.910 ;
        RECT 123.760 158.380 123.930 158.550 ;
        RECT 123.760 158.020 123.930 158.190 ;
        RECT 123.760 157.660 123.930 157.830 ;
        RECT 125.130 159.100 125.300 159.270 ;
        RECT 125.130 158.740 125.300 158.910 ;
        RECT 125.130 158.380 125.300 158.550 ;
        RECT 125.130 158.020 125.300 158.190 ;
        RECT 125.130 157.660 125.300 157.830 ;
        RECT 125.680 158.950 125.850 159.120 ;
        RECT 125.680 158.590 125.850 158.760 ;
        RECT 125.680 158.230 125.850 158.400 ;
        RECT 125.680 157.870 125.850 158.040 ;
        RECT 121.840 157.450 122.010 157.620 ;
        RECT 125.680 157.510 125.850 157.680 ;
        RECT 121.840 157.090 122.010 157.260 ;
        RECT 122.895 157.240 123.065 157.410 ;
        RECT 123.255 157.240 123.425 157.410 ;
        RECT 124.265 157.240 124.435 157.410 ;
        RECT 124.625 157.240 124.795 157.410 ;
        RECT 125.680 157.150 125.850 157.320 ;
        RECT 121.840 156.730 122.010 156.900 ;
        RECT 121.840 156.370 122.010 156.540 ;
        RECT 121.840 156.010 122.010 156.180 ;
        RECT 121.840 155.650 122.010 155.820 ;
        RECT 121.840 155.290 122.010 155.460 ;
        RECT 122.390 156.820 122.560 156.990 ;
        RECT 122.390 156.460 122.560 156.630 ;
        RECT 122.390 156.100 122.560 156.270 ;
        RECT 122.390 155.740 122.560 155.910 ;
        RECT 122.390 155.380 122.560 155.550 ;
        RECT 123.760 156.820 123.930 156.990 ;
        RECT 123.760 156.460 123.930 156.630 ;
        RECT 123.760 156.100 123.930 156.270 ;
        RECT 123.760 155.740 123.930 155.910 ;
        RECT 123.760 155.380 123.930 155.550 ;
        RECT 125.130 156.820 125.300 156.990 ;
        RECT 125.130 156.460 125.300 156.630 ;
        RECT 125.130 156.100 125.300 156.270 ;
        RECT 125.130 155.740 125.300 155.910 ;
        RECT 125.130 155.380 125.300 155.550 ;
        RECT 125.680 156.790 125.850 156.960 ;
        RECT 125.680 156.430 125.850 156.600 ;
        RECT 125.680 156.070 125.850 156.240 ;
        RECT 125.680 155.710 125.850 155.880 ;
        RECT 125.680 155.350 125.850 155.520 ;
        RECT 121.840 154.930 122.010 155.100 ;
        RECT 122.895 154.960 123.065 155.130 ;
        RECT 123.255 154.960 123.425 155.130 ;
        RECT 124.265 154.960 124.435 155.130 ;
        RECT 124.625 154.960 124.795 155.130 ;
        RECT 125.680 154.990 125.850 155.160 ;
        RECT 121.840 154.570 122.010 154.740 ;
        RECT 121.840 154.210 122.010 154.380 ;
        RECT 121.840 153.850 122.010 154.020 ;
        RECT 121.840 153.490 122.010 153.660 ;
        RECT 121.840 153.130 122.010 153.300 ;
        RECT 122.390 154.540 122.560 154.710 ;
        RECT 122.390 154.180 122.560 154.350 ;
        RECT 122.390 153.820 122.560 153.990 ;
        RECT 122.390 153.460 122.560 153.630 ;
        RECT 122.390 153.100 122.560 153.270 ;
        RECT 123.760 154.540 123.930 154.710 ;
        RECT 123.760 154.180 123.930 154.350 ;
        RECT 123.760 153.820 123.930 153.990 ;
        RECT 123.760 153.460 123.930 153.630 ;
        RECT 123.760 153.100 123.930 153.270 ;
        RECT 125.130 154.540 125.300 154.710 ;
        RECT 125.130 154.180 125.300 154.350 ;
        RECT 125.130 153.820 125.300 153.990 ;
        RECT 125.130 153.460 125.300 153.630 ;
        RECT 125.130 153.100 125.300 153.270 ;
        RECT 125.680 154.630 125.850 154.800 ;
        RECT 125.680 154.270 125.850 154.440 ;
        RECT 125.680 153.910 125.850 154.080 ;
        RECT 125.680 153.550 125.850 153.720 ;
        RECT 125.680 153.190 125.850 153.360 ;
        RECT 121.840 152.770 122.010 152.940 ;
        RECT 122.895 152.680 123.065 152.850 ;
        RECT 123.255 152.680 123.425 152.850 ;
        RECT 124.265 152.680 124.435 152.850 ;
        RECT 124.625 152.680 124.795 152.850 ;
        RECT 125.680 152.830 125.850 153.000 ;
        RECT 121.840 152.410 122.010 152.580 ;
        RECT 125.680 152.470 125.850 152.640 ;
        RECT 121.840 152.050 122.010 152.220 ;
        RECT 121.840 151.690 122.010 151.860 ;
        RECT 121.840 151.330 122.010 151.500 ;
        RECT 121.840 150.970 122.010 151.140 ;
        RECT 122.390 152.260 122.560 152.430 ;
        RECT 122.390 151.900 122.560 152.070 ;
        RECT 122.390 151.540 122.560 151.710 ;
        RECT 122.390 151.180 122.560 151.350 ;
        RECT 122.390 150.820 122.560 150.990 ;
        RECT 123.760 152.260 123.930 152.430 ;
        RECT 123.760 151.900 123.930 152.070 ;
        RECT 123.760 151.540 123.930 151.710 ;
        RECT 123.760 151.180 123.930 151.350 ;
        RECT 123.760 150.820 123.930 150.990 ;
        RECT 125.130 152.260 125.300 152.430 ;
        RECT 125.130 151.900 125.300 152.070 ;
        RECT 125.130 151.540 125.300 151.710 ;
        RECT 125.130 151.180 125.300 151.350 ;
        RECT 125.130 150.820 125.300 150.990 ;
        RECT 125.680 152.110 125.850 152.280 ;
        RECT 125.680 151.750 125.850 151.920 ;
        RECT 125.680 151.390 125.850 151.560 ;
        RECT 125.680 151.030 125.850 151.200 ;
        RECT 121.840 150.610 122.010 150.780 ;
        RECT 125.680 150.670 125.850 150.840 ;
        RECT 121.840 150.250 122.010 150.420 ;
        RECT 122.895 150.400 123.065 150.570 ;
        RECT 123.255 150.400 123.425 150.570 ;
        RECT 124.265 150.400 124.435 150.570 ;
        RECT 124.625 150.400 124.795 150.570 ;
        RECT 125.680 150.310 125.850 150.480 ;
        RECT 121.840 149.890 122.010 150.060 ;
        RECT 121.840 149.530 122.010 149.700 ;
        RECT 121.840 149.170 122.010 149.340 ;
        RECT 121.840 148.810 122.010 148.980 ;
        RECT 121.840 148.450 122.010 148.620 ;
        RECT 122.390 149.980 122.560 150.150 ;
        RECT 122.390 149.620 122.560 149.790 ;
        RECT 122.390 149.260 122.560 149.430 ;
        RECT 122.390 148.900 122.560 149.070 ;
        RECT 122.390 148.540 122.560 148.710 ;
        RECT 123.760 149.980 123.930 150.150 ;
        RECT 123.760 149.620 123.930 149.790 ;
        RECT 123.760 149.260 123.930 149.430 ;
        RECT 123.760 148.900 123.930 149.070 ;
        RECT 123.760 148.540 123.930 148.710 ;
        RECT 125.130 149.980 125.300 150.150 ;
        RECT 125.130 149.620 125.300 149.790 ;
        RECT 125.130 149.260 125.300 149.430 ;
        RECT 125.130 148.900 125.300 149.070 ;
        RECT 125.130 148.540 125.300 148.710 ;
        RECT 125.680 149.950 125.850 150.120 ;
        RECT 125.680 149.590 125.850 149.760 ;
        RECT 125.680 149.230 125.850 149.400 ;
        RECT 125.680 148.870 125.850 149.040 ;
        RECT 125.680 148.510 125.850 148.680 ;
        RECT 121.840 148.090 122.010 148.260 ;
        RECT 122.895 148.120 123.065 148.290 ;
        RECT 123.255 148.120 123.425 148.290 ;
        RECT 124.265 148.120 124.435 148.290 ;
        RECT 124.625 148.120 124.795 148.290 ;
        RECT 125.680 148.150 125.850 148.320 ;
        RECT 121.840 147.730 122.010 147.900 ;
        RECT 121.840 147.370 122.010 147.540 ;
        RECT 121.840 147.010 122.010 147.180 ;
        RECT 121.840 146.650 122.010 146.820 ;
        RECT 121.840 146.290 122.010 146.460 ;
        RECT 122.390 147.700 122.560 147.870 ;
        RECT 122.390 147.340 122.560 147.510 ;
        RECT 122.390 146.980 122.560 147.150 ;
        RECT 122.390 146.620 122.560 146.790 ;
        RECT 122.390 146.260 122.560 146.430 ;
        RECT 123.760 147.700 123.930 147.870 ;
        RECT 123.760 147.340 123.930 147.510 ;
        RECT 123.760 146.980 123.930 147.150 ;
        RECT 123.760 146.620 123.930 146.790 ;
        RECT 123.760 146.260 123.930 146.430 ;
        RECT 125.130 147.700 125.300 147.870 ;
        RECT 125.130 147.340 125.300 147.510 ;
        RECT 125.130 146.980 125.300 147.150 ;
        RECT 125.130 146.620 125.300 146.790 ;
        RECT 125.130 146.260 125.300 146.430 ;
        RECT 125.680 147.790 125.850 147.960 ;
        RECT 125.680 147.430 125.850 147.600 ;
        RECT 125.680 147.070 125.850 147.240 ;
        RECT 125.680 146.710 125.850 146.880 ;
        RECT 125.680 146.350 125.850 146.520 ;
        RECT 121.840 145.930 122.010 146.100 ;
        RECT 122.895 145.840 123.065 146.010 ;
        RECT 123.255 145.840 123.425 146.010 ;
        RECT 124.265 145.840 124.435 146.010 ;
        RECT 124.625 145.840 124.795 146.010 ;
        RECT 125.680 145.990 125.850 146.160 ;
        RECT 121.840 145.570 122.010 145.740 ;
        RECT 125.680 145.630 125.850 145.800 ;
        RECT 121.840 145.210 122.010 145.380 ;
        RECT 121.840 144.850 122.010 145.020 ;
        RECT 121.840 144.490 122.010 144.660 ;
        RECT 121.840 144.130 122.010 144.300 ;
        RECT 122.390 145.420 122.560 145.590 ;
        RECT 122.390 145.060 122.560 145.230 ;
        RECT 122.390 144.700 122.560 144.870 ;
        RECT 122.390 144.340 122.560 144.510 ;
        RECT 122.390 143.980 122.560 144.150 ;
        RECT 123.760 145.420 123.930 145.590 ;
        RECT 123.760 145.060 123.930 145.230 ;
        RECT 123.760 144.700 123.930 144.870 ;
        RECT 123.760 144.340 123.930 144.510 ;
        RECT 123.760 143.980 123.930 144.150 ;
        RECT 125.130 145.420 125.300 145.590 ;
        RECT 125.130 145.060 125.300 145.230 ;
        RECT 125.130 144.700 125.300 144.870 ;
        RECT 125.130 144.340 125.300 144.510 ;
        RECT 125.130 143.980 125.300 144.150 ;
        RECT 125.680 145.270 125.850 145.440 ;
        RECT 125.680 144.910 125.850 145.080 ;
        RECT 125.680 144.550 125.850 144.720 ;
        RECT 125.680 144.190 125.850 144.360 ;
        RECT 121.840 143.770 122.010 143.940 ;
        RECT 125.680 143.830 125.850 144.000 ;
        RECT 121.840 143.410 122.010 143.580 ;
        RECT 122.895 143.560 123.065 143.730 ;
        RECT 123.255 143.560 123.425 143.730 ;
        RECT 124.265 143.560 124.435 143.730 ;
        RECT 124.625 143.560 124.795 143.730 ;
        RECT 125.680 143.470 125.850 143.640 ;
        RECT 121.840 143.050 122.010 143.220 ;
        RECT 121.840 142.690 122.010 142.860 ;
        RECT 121.840 142.330 122.010 142.500 ;
        RECT 121.840 141.970 122.010 142.140 ;
        RECT 121.840 141.610 122.010 141.780 ;
        RECT 122.390 143.140 122.560 143.310 ;
        RECT 122.390 142.780 122.560 142.950 ;
        RECT 122.390 142.420 122.560 142.590 ;
        RECT 122.390 142.060 122.560 142.230 ;
        RECT 122.390 141.700 122.560 141.870 ;
        RECT 123.760 143.140 123.930 143.310 ;
        RECT 123.760 142.780 123.930 142.950 ;
        RECT 123.760 142.420 123.930 142.590 ;
        RECT 123.760 142.060 123.930 142.230 ;
        RECT 123.760 141.700 123.930 141.870 ;
        RECT 125.130 143.140 125.300 143.310 ;
        RECT 125.130 142.780 125.300 142.950 ;
        RECT 125.130 142.420 125.300 142.590 ;
        RECT 125.130 142.060 125.300 142.230 ;
        RECT 125.130 141.700 125.300 141.870 ;
        RECT 125.680 143.110 125.850 143.280 ;
        RECT 125.680 142.750 125.850 142.920 ;
        RECT 125.680 142.390 125.850 142.560 ;
        RECT 125.680 142.030 125.850 142.200 ;
        RECT 125.680 141.670 125.850 141.840 ;
        RECT 121.840 141.250 122.010 141.420 ;
        RECT 122.895 141.280 123.065 141.450 ;
        RECT 123.255 141.280 123.425 141.450 ;
        RECT 124.265 141.280 124.435 141.450 ;
        RECT 124.625 141.280 124.795 141.450 ;
        RECT 125.680 141.310 125.850 141.480 ;
        RECT 121.840 140.890 122.010 141.060 ;
        RECT 121.840 140.530 122.010 140.700 ;
        RECT 121.840 140.170 122.010 140.340 ;
        RECT 121.840 139.810 122.010 139.980 ;
        RECT 121.840 139.450 122.010 139.620 ;
        RECT 122.390 140.860 122.560 141.030 ;
        RECT 122.390 140.500 122.560 140.670 ;
        RECT 122.390 140.140 122.560 140.310 ;
        RECT 122.390 139.780 122.560 139.950 ;
        RECT 122.390 139.420 122.560 139.590 ;
        RECT 123.760 140.860 123.930 141.030 ;
        RECT 123.760 140.500 123.930 140.670 ;
        RECT 123.760 140.140 123.930 140.310 ;
        RECT 123.760 139.780 123.930 139.950 ;
        RECT 123.760 139.420 123.930 139.590 ;
        RECT 125.130 140.860 125.300 141.030 ;
        RECT 125.130 140.500 125.300 140.670 ;
        RECT 125.130 140.140 125.300 140.310 ;
        RECT 125.130 139.780 125.300 139.950 ;
        RECT 125.130 139.420 125.300 139.590 ;
        RECT 125.680 140.950 125.850 141.120 ;
        RECT 125.680 140.590 125.850 140.760 ;
        RECT 125.680 140.230 125.850 140.400 ;
        RECT 125.680 139.870 125.850 140.040 ;
        RECT 125.680 139.510 125.850 139.680 ;
        RECT 121.840 139.090 122.010 139.260 ;
        RECT 122.895 139.000 123.065 139.170 ;
        RECT 123.255 139.000 123.425 139.170 ;
        RECT 124.265 139.000 124.435 139.170 ;
        RECT 124.625 139.000 124.795 139.170 ;
        RECT 125.680 139.150 125.850 139.320 ;
        RECT 121.840 138.730 122.010 138.900 ;
        RECT 125.680 138.790 125.850 138.960 ;
        RECT 121.840 138.370 122.010 138.540 ;
        RECT 121.840 138.010 122.010 138.180 ;
        RECT 121.840 137.650 122.010 137.820 ;
        RECT 121.840 137.290 122.010 137.460 ;
        RECT 122.390 138.580 122.560 138.750 ;
        RECT 122.390 138.220 122.560 138.390 ;
        RECT 122.390 137.860 122.560 138.030 ;
        RECT 122.390 137.500 122.560 137.670 ;
        RECT 122.390 137.140 122.560 137.310 ;
        RECT 123.760 138.580 123.930 138.750 ;
        RECT 123.760 138.220 123.930 138.390 ;
        RECT 123.760 137.860 123.930 138.030 ;
        RECT 123.760 137.500 123.930 137.670 ;
        RECT 123.760 137.140 123.930 137.310 ;
        RECT 125.130 138.580 125.300 138.750 ;
        RECT 125.130 138.220 125.300 138.390 ;
        RECT 125.130 137.860 125.300 138.030 ;
        RECT 125.130 137.500 125.300 137.670 ;
        RECT 125.130 137.140 125.300 137.310 ;
        RECT 125.680 138.430 125.850 138.600 ;
        RECT 125.680 138.070 125.850 138.240 ;
        RECT 125.680 137.710 125.850 137.880 ;
        RECT 125.680 137.350 125.850 137.520 ;
        RECT 121.840 136.930 122.010 137.100 ;
        RECT 125.680 136.990 125.850 137.160 ;
        RECT 121.840 136.570 122.010 136.740 ;
        RECT 122.895 136.720 123.065 136.890 ;
        RECT 123.255 136.720 123.425 136.890 ;
        RECT 124.265 136.720 124.435 136.890 ;
        RECT 124.625 136.720 124.795 136.890 ;
        RECT 125.680 136.630 125.850 136.800 ;
        RECT 121.840 136.210 122.010 136.380 ;
        RECT 121.840 135.850 122.010 136.020 ;
        RECT 121.840 135.490 122.010 135.660 ;
        RECT 121.840 135.130 122.010 135.300 ;
        RECT 121.840 134.770 122.010 134.940 ;
        RECT 122.390 136.300 122.560 136.470 ;
        RECT 122.390 135.940 122.560 136.110 ;
        RECT 122.390 135.580 122.560 135.750 ;
        RECT 122.390 135.220 122.560 135.390 ;
        RECT 122.390 134.860 122.560 135.030 ;
        RECT 123.760 136.300 123.930 136.470 ;
        RECT 123.760 135.940 123.930 136.110 ;
        RECT 123.760 135.580 123.930 135.750 ;
        RECT 123.760 135.220 123.930 135.390 ;
        RECT 123.760 134.860 123.930 135.030 ;
        RECT 125.130 136.300 125.300 136.470 ;
        RECT 125.130 135.940 125.300 136.110 ;
        RECT 125.130 135.580 125.300 135.750 ;
        RECT 125.130 135.220 125.300 135.390 ;
        RECT 125.130 134.860 125.300 135.030 ;
        RECT 125.680 136.270 125.850 136.440 ;
        RECT 125.680 135.910 125.850 136.080 ;
        RECT 125.680 135.550 125.850 135.720 ;
        RECT 125.680 135.190 125.850 135.360 ;
        RECT 125.680 134.830 125.850 135.000 ;
        RECT 121.840 134.410 122.010 134.580 ;
        RECT 122.895 134.440 123.065 134.610 ;
        RECT 123.255 134.440 123.425 134.610 ;
        RECT 124.265 134.440 124.435 134.610 ;
        RECT 124.625 134.440 124.795 134.610 ;
        RECT 125.680 134.470 125.850 134.640 ;
        RECT 121.840 134.050 122.010 134.220 ;
        RECT 121.840 133.690 122.010 133.860 ;
        RECT 121.840 133.330 122.010 133.500 ;
        RECT 121.840 132.970 122.010 133.140 ;
        RECT 121.840 132.610 122.010 132.780 ;
        RECT 122.390 134.020 122.560 134.190 ;
        RECT 122.390 133.660 122.560 133.830 ;
        RECT 122.390 133.300 122.560 133.470 ;
        RECT 122.390 132.940 122.560 133.110 ;
        RECT 122.390 132.580 122.560 132.750 ;
        RECT 123.760 134.020 123.930 134.190 ;
        RECT 123.760 133.660 123.930 133.830 ;
        RECT 123.760 133.300 123.930 133.470 ;
        RECT 123.760 132.940 123.930 133.110 ;
        RECT 123.760 132.580 123.930 132.750 ;
        RECT 125.130 134.020 125.300 134.190 ;
        RECT 125.130 133.660 125.300 133.830 ;
        RECT 125.130 133.300 125.300 133.470 ;
        RECT 125.130 132.940 125.300 133.110 ;
        RECT 125.130 132.580 125.300 132.750 ;
        RECT 125.680 134.110 125.850 134.280 ;
        RECT 125.680 133.750 125.850 133.920 ;
        RECT 125.680 133.390 125.850 133.560 ;
        RECT 125.680 133.030 125.850 133.200 ;
        RECT 125.680 132.670 125.850 132.840 ;
        RECT 121.840 132.250 122.010 132.420 ;
        RECT 122.895 132.160 123.065 132.330 ;
        RECT 123.255 132.160 123.425 132.330 ;
        RECT 124.265 132.160 124.435 132.330 ;
        RECT 124.625 132.160 124.795 132.330 ;
        RECT 125.680 132.310 125.850 132.480 ;
        RECT 121.840 131.890 122.010 132.060 ;
        RECT 125.680 131.950 125.850 132.120 ;
        RECT 121.840 131.530 122.010 131.700 ;
        RECT 121.840 131.170 122.010 131.340 ;
        RECT 121.840 130.810 122.010 130.980 ;
        RECT 121.840 130.450 122.010 130.620 ;
        RECT 122.390 131.740 122.560 131.910 ;
        RECT 122.390 131.380 122.560 131.550 ;
        RECT 122.390 131.020 122.560 131.190 ;
        RECT 122.390 130.660 122.560 130.830 ;
        RECT 122.390 130.300 122.560 130.470 ;
        RECT 123.760 131.740 123.930 131.910 ;
        RECT 123.760 131.380 123.930 131.550 ;
        RECT 123.760 131.020 123.930 131.190 ;
        RECT 123.760 130.660 123.930 130.830 ;
        RECT 123.760 130.300 123.930 130.470 ;
        RECT 125.130 131.740 125.300 131.910 ;
        RECT 125.130 131.380 125.300 131.550 ;
        RECT 125.130 131.020 125.300 131.190 ;
        RECT 125.130 130.660 125.300 130.830 ;
        RECT 125.130 130.300 125.300 130.470 ;
        RECT 125.680 131.590 125.850 131.760 ;
        RECT 125.680 131.230 125.850 131.400 ;
        RECT 125.680 130.870 125.850 131.040 ;
        RECT 125.680 130.510 125.850 130.680 ;
        RECT 121.840 130.090 122.010 130.260 ;
        RECT 125.680 130.150 125.850 130.320 ;
        RECT 121.840 129.730 122.010 129.900 ;
        RECT 122.895 129.880 123.065 130.050 ;
        RECT 123.255 129.880 123.425 130.050 ;
        RECT 124.265 129.880 124.435 130.050 ;
        RECT 124.625 129.880 124.795 130.050 ;
        RECT 125.680 129.790 125.850 129.960 ;
        RECT 121.840 129.370 122.010 129.540 ;
        RECT 121.840 129.010 122.010 129.180 ;
        RECT 121.840 128.650 122.010 128.820 ;
        RECT 121.840 128.290 122.010 128.460 ;
        RECT 121.840 127.930 122.010 128.100 ;
        RECT 122.390 129.460 122.560 129.630 ;
        RECT 122.390 129.100 122.560 129.270 ;
        RECT 122.390 128.740 122.560 128.910 ;
        RECT 122.390 128.380 122.560 128.550 ;
        RECT 122.390 128.020 122.560 128.190 ;
        RECT 123.760 129.460 123.930 129.630 ;
        RECT 123.760 129.100 123.930 129.270 ;
        RECT 123.760 128.740 123.930 128.910 ;
        RECT 123.760 128.380 123.930 128.550 ;
        RECT 123.760 128.020 123.930 128.190 ;
        RECT 125.130 129.460 125.300 129.630 ;
        RECT 125.130 129.100 125.300 129.270 ;
        RECT 125.130 128.740 125.300 128.910 ;
        RECT 125.130 128.380 125.300 128.550 ;
        RECT 125.130 128.020 125.300 128.190 ;
        RECT 125.680 129.430 125.850 129.600 ;
        RECT 125.680 129.070 125.850 129.240 ;
        RECT 125.680 128.710 125.850 128.880 ;
        RECT 125.680 128.350 125.850 128.520 ;
        RECT 125.680 127.990 125.850 128.160 ;
        RECT 121.840 127.570 122.010 127.740 ;
        RECT 122.895 127.600 123.065 127.770 ;
        RECT 123.255 127.600 123.425 127.770 ;
        RECT 124.265 127.600 124.435 127.770 ;
        RECT 124.625 127.600 124.795 127.770 ;
        RECT 125.680 127.630 125.850 127.800 ;
        RECT 121.840 127.210 122.010 127.380 ;
        RECT 121.840 126.850 122.010 127.020 ;
        RECT 121.840 126.490 122.010 126.660 ;
        RECT 121.840 126.130 122.010 126.300 ;
        RECT 121.840 125.770 122.010 125.940 ;
        RECT 122.390 127.180 122.560 127.350 ;
        RECT 122.390 126.820 122.560 126.990 ;
        RECT 122.390 126.460 122.560 126.630 ;
        RECT 122.390 126.100 122.560 126.270 ;
        RECT 122.390 125.740 122.560 125.910 ;
        RECT 123.760 127.180 123.930 127.350 ;
        RECT 123.760 126.820 123.930 126.990 ;
        RECT 123.760 126.460 123.930 126.630 ;
        RECT 123.760 126.100 123.930 126.270 ;
        RECT 123.760 125.740 123.930 125.910 ;
        RECT 125.130 127.180 125.300 127.350 ;
        RECT 125.130 126.820 125.300 126.990 ;
        RECT 125.130 126.460 125.300 126.630 ;
        RECT 125.130 126.100 125.300 126.270 ;
        RECT 125.130 125.740 125.300 125.910 ;
        RECT 125.680 127.270 125.850 127.440 ;
        RECT 125.680 126.910 125.850 127.080 ;
        RECT 125.680 126.550 125.850 126.720 ;
        RECT 125.680 126.190 125.850 126.360 ;
        RECT 125.680 125.830 125.850 126.000 ;
        RECT 121.840 125.410 122.010 125.580 ;
        RECT 122.895 125.320 123.065 125.490 ;
        RECT 123.255 125.320 123.425 125.490 ;
        RECT 124.265 125.320 124.435 125.490 ;
        RECT 124.625 125.320 124.795 125.490 ;
        RECT 125.680 125.470 125.850 125.640 ;
        RECT 121.840 125.050 122.010 125.220 ;
        RECT 125.680 125.110 125.850 125.280 ;
        RECT 121.840 124.690 122.010 124.860 ;
        RECT 121.840 124.330 122.010 124.500 ;
        RECT 121.840 123.970 122.010 124.140 ;
        RECT 121.840 123.610 122.010 123.780 ;
        RECT 122.390 124.900 122.560 125.070 ;
        RECT 122.390 124.540 122.560 124.710 ;
        RECT 122.390 124.180 122.560 124.350 ;
        RECT 122.390 123.820 122.560 123.990 ;
        RECT 122.390 123.460 122.560 123.630 ;
        RECT 123.760 124.900 123.930 125.070 ;
        RECT 123.760 124.540 123.930 124.710 ;
        RECT 123.760 124.180 123.930 124.350 ;
        RECT 123.760 123.820 123.930 123.990 ;
        RECT 123.760 123.460 123.930 123.630 ;
        RECT 125.130 124.900 125.300 125.070 ;
        RECT 125.130 124.540 125.300 124.710 ;
        RECT 125.130 124.180 125.300 124.350 ;
        RECT 125.130 123.820 125.300 123.990 ;
        RECT 125.130 123.460 125.300 123.630 ;
        RECT 125.680 124.750 125.850 124.920 ;
        RECT 125.680 124.390 125.850 124.560 ;
        RECT 125.680 124.030 125.850 124.200 ;
        RECT 125.680 123.670 125.850 123.840 ;
        RECT 121.840 123.250 122.010 123.420 ;
        RECT 125.680 123.310 125.850 123.480 ;
        RECT 121.840 122.890 122.010 123.060 ;
        RECT 122.895 123.040 123.065 123.210 ;
        RECT 123.255 123.040 123.425 123.210 ;
        RECT 124.265 123.040 124.435 123.210 ;
        RECT 124.625 123.040 124.795 123.210 ;
        RECT 125.680 122.950 125.850 123.120 ;
        RECT 121.840 122.530 122.010 122.700 ;
        RECT 121.840 122.170 122.010 122.340 ;
        RECT 121.840 121.810 122.010 121.980 ;
        RECT 121.840 121.450 122.010 121.620 ;
        RECT 121.840 121.090 122.010 121.260 ;
        RECT 122.390 122.620 122.560 122.790 ;
        RECT 122.390 122.260 122.560 122.430 ;
        RECT 122.390 121.900 122.560 122.070 ;
        RECT 122.390 121.540 122.560 121.710 ;
        RECT 122.390 121.180 122.560 121.350 ;
        RECT 123.760 122.620 123.930 122.790 ;
        RECT 123.760 122.260 123.930 122.430 ;
        RECT 123.760 121.900 123.930 122.070 ;
        RECT 123.760 121.540 123.930 121.710 ;
        RECT 123.760 121.180 123.930 121.350 ;
        RECT 125.130 122.620 125.300 122.790 ;
        RECT 125.130 122.260 125.300 122.430 ;
        RECT 125.130 121.900 125.300 122.070 ;
        RECT 125.130 121.540 125.300 121.710 ;
        RECT 125.130 121.180 125.300 121.350 ;
        RECT 125.680 122.590 125.850 122.760 ;
        RECT 125.680 122.230 125.850 122.400 ;
        RECT 125.680 121.870 125.850 122.040 ;
        RECT 125.680 121.510 125.850 121.680 ;
        RECT 125.680 121.150 125.850 121.320 ;
        RECT 122.895 120.760 123.065 120.930 ;
        RECT 123.255 120.760 123.425 120.930 ;
        RECT 124.265 120.760 124.435 120.930 ;
        RECT 124.625 120.760 124.795 120.930 ;
        RECT 125.680 120.790 125.850 120.960 ;
        RECT 121.840 120.580 122.010 120.750 ;
        RECT 121.840 120.220 122.010 120.390 ;
        RECT 121.840 119.860 122.010 120.030 ;
        RECT 121.840 119.500 122.010 119.670 ;
        RECT 121.840 119.140 122.010 119.310 ;
        RECT 121.840 118.780 122.010 118.950 ;
        RECT 122.390 120.340 122.560 120.510 ;
        RECT 122.390 119.980 122.560 120.150 ;
        RECT 122.390 119.620 122.560 119.790 ;
        RECT 122.390 119.260 122.560 119.430 ;
        RECT 122.390 118.900 122.560 119.070 ;
        RECT 123.760 120.340 123.930 120.510 ;
        RECT 123.760 119.980 123.930 120.150 ;
        RECT 123.760 119.620 123.930 119.790 ;
        RECT 123.760 119.260 123.930 119.430 ;
        RECT 123.760 118.900 123.930 119.070 ;
        RECT 125.130 120.340 125.300 120.510 ;
        RECT 125.130 119.980 125.300 120.150 ;
        RECT 125.130 119.620 125.300 119.790 ;
        RECT 125.130 119.260 125.300 119.430 ;
        RECT 125.130 118.900 125.300 119.070 ;
        RECT 125.680 120.430 125.850 120.600 ;
        RECT 125.680 120.070 125.850 120.240 ;
        RECT 125.680 119.710 125.850 119.880 ;
        RECT 125.680 119.350 125.850 119.520 ;
        RECT 125.680 118.990 125.850 119.160 ;
        RECT 121.840 118.420 122.010 118.590 ;
        RECT 122.895 118.480 123.065 118.650 ;
        RECT 123.255 118.480 123.425 118.650 ;
        RECT 124.265 118.480 124.435 118.650 ;
        RECT 124.625 118.480 124.795 118.650 ;
        RECT 125.680 118.630 125.850 118.800 ;
        RECT 108.635 117.890 108.805 118.060 ;
        RECT 108.635 117.530 108.805 117.700 ;
        RECT 108.635 117.170 108.805 117.340 ;
        RECT 108.635 116.810 108.805 116.980 ;
        RECT 110.555 118.060 110.725 118.230 ;
        RECT 110.555 117.700 110.725 117.870 ;
        RECT 110.555 117.340 110.725 117.510 ;
        RECT 110.555 116.980 110.725 117.150 ;
        RECT 110.555 116.620 110.725 116.790 ;
        RECT 111.925 118.060 112.095 118.230 ;
        RECT 111.925 117.700 112.095 117.870 ;
        RECT 111.925 117.340 112.095 117.510 ;
        RECT 111.925 116.980 112.095 117.150 ;
        RECT 111.925 116.620 112.095 116.790 ;
        RECT 113.845 117.870 114.015 118.040 ;
        RECT 113.845 117.510 114.015 117.680 ;
        RECT 113.845 117.150 114.015 117.320 ;
        RECT 113.845 116.790 114.015 116.960 ;
        RECT 108.635 116.450 108.805 116.620 ;
        RECT 113.845 116.430 114.015 116.600 ;
        RECT 108.635 116.090 108.805 116.260 ;
        RECT 109.690 116.200 109.860 116.370 ;
        RECT 110.050 116.200 110.220 116.370 ;
        RECT 111.060 116.200 111.230 116.370 ;
        RECT 111.420 116.200 111.590 116.370 ;
        RECT 112.430 116.200 112.600 116.370 ;
        RECT 112.790 116.200 112.960 116.370 ;
        RECT 113.845 116.070 114.015 116.240 ;
        RECT 108.635 115.730 108.805 115.900 ;
        RECT 108.635 115.370 108.805 115.540 ;
        RECT 108.635 115.010 108.805 115.180 ;
        RECT 108.635 114.650 108.805 114.820 ;
        RECT 108.635 114.290 108.805 114.460 ;
        RECT 110.555 115.780 110.725 115.950 ;
        RECT 110.555 115.420 110.725 115.590 ;
        RECT 110.555 115.060 110.725 115.230 ;
        RECT 110.555 114.700 110.725 114.870 ;
        RECT 110.555 114.340 110.725 114.510 ;
        RECT 111.925 115.780 112.095 115.950 ;
        RECT 111.925 115.420 112.095 115.590 ;
        RECT 111.925 115.060 112.095 115.230 ;
        RECT 111.925 114.700 112.095 114.870 ;
        RECT 111.925 114.340 112.095 114.510 ;
        RECT 113.845 115.710 114.015 115.880 ;
        RECT 113.845 115.350 114.015 115.520 ;
        RECT 113.845 114.990 114.015 115.160 ;
        RECT 113.845 114.630 114.015 114.800 ;
        RECT 113.845 114.270 114.015 114.440 ;
        RECT 114.925 118.095 115.095 118.265 ;
        RECT 115.535 118.155 115.705 118.325 ;
        RECT 115.895 118.155 116.065 118.325 ;
        RECT 116.255 118.155 116.425 118.325 ;
        RECT 116.615 118.155 116.785 118.325 ;
        RECT 116.975 118.155 117.145 118.325 ;
        RECT 117.335 118.155 117.505 118.325 ;
        RECT 114.925 117.735 115.095 117.905 ;
        RECT 125.680 118.270 125.850 118.440 ;
        RECT 114.925 117.375 115.095 117.545 ;
        RECT 115.980 117.525 116.150 117.695 ;
        RECT 116.340 117.525 116.510 117.695 ;
        RECT 117.395 117.615 117.565 117.785 ;
        RECT 114.925 117.015 115.095 117.185 ;
        RECT 115.980 117.095 116.150 117.265 ;
        RECT 116.340 117.095 116.510 117.265 ;
        RECT 116.845 117.095 117.015 117.265 ;
        RECT 117.395 117.255 117.565 117.425 ;
        RECT 117.395 116.895 117.565 117.065 ;
        RECT 114.925 116.655 115.095 116.825 ;
        RECT 115.980 116.665 116.150 116.835 ;
        RECT 116.340 116.665 116.510 116.835 ;
        RECT 117.395 116.535 117.565 116.705 ;
        RECT 115.475 116.235 115.645 116.405 ;
        RECT 115.980 116.235 116.150 116.405 ;
        RECT 116.340 116.235 116.510 116.405 ;
        RECT 114.925 116.055 115.095 116.225 ;
        RECT 117.395 116.175 117.565 116.345 ;
        RECT 114.925 115.695 115.095 115.865 ;
        RECT 115.980 115.805 116.150 115.975 ;
        RECT 116.340 115.805 116.510 115.975 ;
        RECT 117.395 115.815 117.565 115.985 ;
        RECT 114.925 115.335 115.095 115.505 ;
        RECT 115.980 115.375 116.150 115.545 ;
        RECT 116.340 115.375 116.510 115.545 ;
        RECT 116.845 115.375 117.015 115.545 ;
        RECT 117.395 115.455 117.565 115.625 ;
        RECT 114.925 114.975 115.095 115.145 ;
        RECT 115.980 114.945 116.150 115.115 ;
        RECT 116.340 114.945 116.510 115.115 ;
        RECT 117.395 115.095 117.565 115.265 ;
        RECT 117.395 114.735 117.565 114.905 ;
        RECT 114.985 114.315 115.155 114.485 ;
        RECT 115.345 114.315 115.515 114.485 ;
        RECT 115.705 114.315 115.875 114.485 ;
        RECT 116.065 114.315 116.235 114.485 ;
        RECT 116.425 114.315 116.595 114.485 ;
        RECT 116.785 114.315 116.955 114.485 ;
        RECT 117.395 114.375 117.565 114.545 ;
        RECT 118.195 117.860 118.365 118.030 ;
        RECT 118.745 117.920 118.915 118.090 ;
        RECT 119.105 117.920 119.275 118.090 ;
        RECT 119.465 117.920 119.635 118.090 ;
        RECT 119.825 117.920 119.995 118.090 ;
        RECT 120.185 117.920 120.355 118.090 ;
        RECT 120.545 117.920 120.715 118.090 ;
        RECT 120.905 117.920 121.075 118.090 ;
        RECT 118.195 117.500 118.365 117.670 ;
        RECT 118.195 117.140 118.365 117.310 ;
        RECT 119.400 117.290 119.570 117.460 ;
        RECT 119.760 117.290 119.930 117.460 ;
        RECT 120.965 117.400 121.135 117.570 ;
        RECT 120.965 117.040 121.135 117.210 ;
        RECT 118.195 116.780 118.365 116.950 ;
        RECT 118.745 116.860 118.915 117.030 ;
        RECT 119.400 116.860 119.570 117.030 ;
        RECT 119.760 116.860 119.930 117.030 ;
        RECT 120.965 116.680 121.135 116.850 ;
        RECT 118.195 116.420 118.365 116.590 ;
        RECT 119.400 116.430 119.570 116.600 ;
        RECT 119.760 116.430 119.930 116.600 ;
        RECT 118.195 116.060 118.365 116.230 ;
        RECT 120.965 116.320 121.135 116.490 ;
        RECT 118.745 116.000 118.915 116.170 ;
        RECT 119.400 116.000 119.570 116.170 ;
        RECT 119.760 116.000 119.930 116.170 ;
        RECT 118.195 115.700 118.365 115.870 ;
        RECT 120.965 115.960 121.135 116.130 ;
        RECT 119.400 115.570 119.570 115.740 ;
        RECT 119.760 115.570 119.930 115.740 ;
        RECT 120.965 115.600 121.135 115.770 ;
        RECT 118.195 115.340 118.365 115.510 ;
        RECT 118.195 114.980 118.365 115.150 ;
        RECT 118.745 115.140 118.915 115.310 ;
        RECT 119.400 115.140 119.570 115.310 ;
        RECT 119.760 115.140 119.930 115.310 ;
        RECT 120.965 115.240 121.135 115.410 ;
        RECT 120.965 114.880 121.135 115.050 ;
        RECT 118.195 114.620 118.365 114.790 ;
        RECT 119.400 114.710 119.570 114.880 ;
        RECT 119.760 114.710 119.930 114.880 ;
        RECT 120.965 114.520 121.135 114.690 ;
        RECT 109.690 113.920 109.860 114.090 ;
        RECT 110.050 113.920 110.220 114.090 ;
        RECT 111.060 113.920 111.230 114.090 ;
        RECT 111.420 113.920 111.590 114.090 ;
        RECT 112.430 113.920 112.600 114.090 ;
        RECT 112.790 113.920 112.960 114.090 ;
        RECT 108.635 113.740 108.805 113.910 ;
        RECT 113.845 113.910 114.015 114.080 ;
        RECT 108.635 113.380 108.805 113.550 ;
        RECT 108.635 113.020 108.805 113.190 ;
        RECT 108.635 112.660 108.805 112.830 ;
        RECT 108.635 112.300 108.805 112.470 ;
        RECT 94.935 111.550 95.105 111.720 ;
        RECT 94.935 111.190 95.105 111.360 ;
        RECT 94.935 110.830 95.105 111.000 ;
        RECT 88.545 110.470 88.715 110.640 ;
        RECT 89.340 110.390 89.510 110.560 ;
        RECT 93.710 110.390 93.880 110.560 ;
        RECT 94.070 110.390 94.240 110.560 ;
        RECT 94.935 110.470 95.105 110.640 ;
        RECT 88.545 110.110 88.715 110.280 ;
        RECT 88.545 109.750 88.715 109.920 ;
        RECT 88.545 109.390 88.715 109.560 ;
        RECT 88.545 109.030 88.715 109.200 ;
        RECT 88.545 108.670 88.715 108.840 ;
        RECT 89.925 109.970 90.095 110.140 ;
        RECT 89.925 109.610 90.095 109.780 ;
        RECT 89.925 109.250 90.095 109.420 ;
        RECT 89.925 108.890 90.095 109.060 ;
        RECT 89.925 108.530 90.095 108.700 ;
        RECT 93.055 109.970 93.225 110.140 ;
        RECT 93.055 109.610 93.225 109.780 ;
        RECT 93.055 109.250 93.225 109.420 ;
        RECT 93.055 108.890 93.225 109.060 ;
        RECT 93.055 108.530 93.225 108.700 ;
        RECT 94.935 110.110 95.105 110.280 ;
        RECT 94.935 109.750 95.105 109.920 ;
        RECT 94.935 109.390 95.105 109.560 ;
        RECT 94.935 109.030 95.105 109.200 ;
        RECT 94.935 108.670 95.105 108.840 ;
        RECT 88.545 108.310 88.715 108.480 ;
        RECT 94.935 108.310 95.105 108.480 ;
        RECT 88.545 107.950 88.715 108.120 ;
        RECT 89.340 108.110 89.510 108.280 ;
        RECT 93.710 108.110 93.880 108.280 ;
        RECT 94.070 108.110 94.240 108.280 ;
        RECT 94.935 107.950 95.105 108.120 ;
        RECT 88.545 107.590 88.715 107.760 ;
        RECT 88.545 107.230 88.715 107.400 ;
        RECT 88.545 106.870 88.715 107.040 ;
        RECT 88.545 106.510 88.715 106.680 ;
        RECT 88.545 106.150 88.715 106.320 ;
        RECT 89.925 107.690 90.095 107.860 ;
        RECT 89.925 107.330 90.095 107.500 ;
        RECT 89.925 106.970 90.095 107.140 ;
        RECT 89.925 106.610 90.095 106.780 ;
        RECT 89.925 106.250 90.095 106.420 ;
        RECT 93.055 107.690 93.225 107.860 ;
        RECT 93.055 107.330 93.225 107.500 ;
        RECT 93.055 106.970 93.225 107.140 ;
        RECT 93.055 106.610 93.225 106.780 ;
        RECT 93.055 106.250 93.225 106.420 ;
        RECT 94.935 107.590 95.105 107.760 ;
        RECT 94.935 107.230 95.105 107.400 ;
        RECT 94.935 106.870 95.105 107.040 ;
        RECT 94.935 106.510 95.105 106.680 ;
        RECT 94.935 106.150 95.105 106.320 ;
        RECT 88.545 105.790 88.715 105.960 ;
        RECT 89.340 105.830 89.510 106.000 ;
        RECT 93.710 105.830 93.880 106.000 ;
        RECT 94.070 105.830 94.240 106.000 ;
        RECT 88.545 105.430 88.715 105.600 ;
        RECT 94.935 105.790 95.105 105.960 ;
        RECT 88.545 105.070 88.715 105.240 ;
        RECT 88.545 104.710 88.715 104.880 ;
        RECT 88.545 104.350 88.715 104.520 ;
        RECT 88.545 103.990 88.715 104.160 ;
        RECT 89.925 105.410 90.095 105.580 ;
        RECT 89.925 105.050 90.095 105.220 ;
        RECT 89.925 104.690 90.095 104.860 ;
        RECT 89.925 104.330 90.095 104.500 ;
        RECT 89.925 103.970 90.095 104.140 ;
        RECT 93.055 105.410 93.225 105.580 ;
        RECT 93.055 105.050 93.225 105.220 ;
        RECT 93.055 104.690 93.225 104.860 ;
        RECT 93.055 104.330 93.225 104.500 ;
        RECT 93.055 103.970 93.225 104.140 ;
        RECT 94.935 105.430 95.105 105.600 ;
        RECT 94.935 105.070 95.105 105.240 ;
        RECT 94.935 104.710 95.105 104.880 ;
        RECT 94.935 104.350 95.105 104.520 ;
        RECT 94.935 103.990 95.105 104.160 ;
        RECT 88.545 103.630 88.715 103.800 ;
        RECT 89.340 103.550 89.510 103.720 ;
        RECT 93.710 103.550 93.880 103.720 ;
        RECT 94.070 103.550 94.240 103.720 ;
        RECT 94.935 103.630 95.105 103.800 ;
        RECT 88.545 103.270 88.715 103.440 ;
        RECT 88.545 102.910 88.715 103.080 ;
        RECT 88.545 102.550 88.715 102.720 ;
        RECT 88.545 102.190 88.715 102.360 ;
        RECT 88.545 101.830 88.715 102.000 ;
        RECT 89.925 103.130 90.095 103.300 ;
        RECT 89.925 102.770 90.095 102.940 ;
        RECT 89.925 102.410 90.095 102.580 ;
        RECT 89.925 102.050 90.095 102.220 ;
        RECT 89.925 101.690 90.095 101.860 ;
        RECT 93.055 103.130 93.225 103.300 ;
        RECT 93.055 102.770 93.225 102.940 ;
        RECT 93.055 102.410 93.225 102.580 ;
        RECT 93.055 102.050 93.225 102.220 ;
        RECT 93.055 101.690 93.225 101.860 ;
        RECT 94.935 103.270 95.105 103.440 ;
        RECT 94.935 102.910 95.105 103.080 ;
        RECT 94.935 102.550 95.105 102.720 ;
        RECT 94.935 102.190 95.105 102.360 ;
        RECT 94.935 101.830 95.105 102.000 ;
        RECT 88.545 101.470 88.715 101.640 ;
        RECT 94.935 101.470 95.105 101.640 ;
        RECT 88.545 101.110 88.715 101.280 ;
        RECT 89.340 101.270 89.510 101.440 ;
        RECT 93.710 101.270 93.880 101.440 ;
        RECT 94.070 101.270 94.240 101.440 ;
        RECT 94.935 101.110 95.105 101.280 ;
        RECT 88.545 100.750 88.715 100.920 ;
        RECT 88.545 100.390 88.715 100.560 ;
        RECT 88.545 100.030 88.715 100.200 ;
        RECT 88.545 99.670 88.715 99.840 ;
        RECT 88.545 99.310 88.715 99.480 ;
        RECT 89.925 100.850 90.095 101.020 ;
        RECT 89.925 100.490 90.095 100.660 ;
        RECT 89.925 100.130 90.095 100.300 ;
        RECT 89.925 99.770 90.095 99.940 ;
        RECT 89.925 99.410 90.095 99.580 ;
        RECT 93.055 100.850 93.225 101.020 ;
        RECT 93.055 100.490 93.225 100.660 ;
        RECT 93.055 100.130 93.225 100.300 ;
        RECT 93.055 99.770 93.225 99.940 ;
        RECT 93.055 99.410 93.225 99.580 ;
        RECT 94.935 100.750 95.105 100.920 ;
        RECT 94.935 100.390 95.105 100.560 ;
        RECT 94.935 100.030 95.105 100.200 ;
        RECT 94.935 99.670 95.105 99.840 ;
        RECT 94.935 99.310 95.105 99.480 ;
        RECT 88.545 98.950 88.715 99.120 ;
        RECT 89.340 98.990 89.510 99.160 ;
        RECT 93.710 98.990 93.880 99.160 ;
        RECT 94.070 98.990 94.240 99.160 ;
        RECT 88.545 98.590 88.715 98.760 ;
        RECT 94.935 98.950 95.105 99.120 ;
        RECT 88.545 98.230 88.715 98.400 ;
        RECT 88.545 97.870 88.715 98.040 ;
        RECT 88.545 97.510 88.715 97.680 ;
        RECT 88.545 97.150 88.715 97.320 ;
        RECT 89.925 98.570 90.095 98.740 ;
        RECT 89.925 98.210 90.095 98.380 ;
        RECT 89.925 97.850 90.095 98.020 ;
        RECT 89.925 97.490 90.095 97.660 ;
        RECT 89.925 97.130 90.095 97.300 ;
        RECT 93.055 98.570 93.225 98.740 ;
        RECT 93.055 98.210 93.225 98.380 ;
        RECT 93.055 97.850 93.225 98.020 ;
        RECT 93.055 97.490 93.225 97.660 ;
        RECT 93.055 97.130 93.225 97.300 ;
        RECT 94.935 98.590 95.105 98.760 ;
        RECT 94.935 98.230 95.105 98.400 ;
        RECT 94.935 97.870 95.105 98.040 ;
        RECT 94.935 97.510 95.105 97.680 ;
        RECT 94.935 97.150 95.105 97.320 ;
        RECT 88.545 96.790 88.715 96.960 ;
        RECT 89.340 96.710 89.510 96.880 ;
        RECT 93.710 96.710 93.880 96.880 ;
        RECT 94.070 96.710 94.240 96.880 ;
        RECT 94.935 96.790 95.105 96.960 ;
        RECT 88.545 96.430 88.715 96.600 ;
        RECT 88.545 96.070 88.715 96.240 ;
        RECT 88.545 95.710 88.715 95.880 ;
        RECT 88.545 95.350 88.715 95.520 ;
        RECT 88.545 94.990 88.715 95.160 ;
        RECT 89.925 96.290 90.095 96.460 ;
        RECT 89.925 95.930 90.095 96.100 ;
        RECT 89.925 95.570 90.095 95.740 ;
        RECT 89.925 95.210 90.095 95.380 ;
        RECT 89.925 94.850 90.095 95.020 ;
        RECT 93.055 96.290 93.225 96.460 ;
        RECT 93.055 95.930 93.225 96.100 ;
        RECT 93.055 95.570 93.225 95.740 ;
        RECT 93.055 95.210 93.225 95.380 ;
        RECT 93.055 94.850 93.225 95.020 ;
        RECT 94.935 96.430 95.105 96.600 ;
        RECT 94.935 96.070 95.105 96.240 ;
        RECT 94.935 95.710 95.105 95.880 ;
        RECT 94.935 95.350 95.105 95.520 ;
        RECT 94.935 94.990 95.105 95.160 ;
        RECT 88.545 94.630 88.715 94.800 ;
        RECT 94.935 94.630 95.105 94.800 ;
        RECT 88.545 94.270 88.715 94.440 ;
        RECT 89.340 94.430 89.510 94.600 ;
        RECT 93.710 94.430 93.880 94.600 ;
        RECT 94.070 94.430 94.240 94.600 ;
        RECT 94.935 94.270 95.105 94.440 ;
        RECT 88.545 93.910 88.715 94.080 ;
        RECT 88.545 93.550 88.715 93.720 ;
        RECT 88.545 93.190 88.715 93.360 ;
        RECT 88.545 92.830 88.715 93.000 ;
        RECT 88.545 92.470 88.715 92.640 ;
        RECT 89.925 94.010 90.095 94.180 ;
        RECT 89.925 93.650 90.095 93.820 ;
        RECT 89.925 93.290 90.095 93.460 ;
        RECT 89.925 92.930 90.095 93.100 ;
        RECT 89.925 92.570 90.095 92.740 ;
        RECT 93.055 94.010 93.225 94.180 ;
        RECT 93.055 93.650 93.225 93.820 ;
        RECT 93.055 93.290 93.225 93.460 ;
        RECT 93.055 92.930 93.225 93.100 ;
        RECT 93.055 92.570 93.225 92.740 ;
        RECT 94.935 93.910 95.105 94.080 ;
        RECT 94.935 93.550 95.105 93.720 ;
        RECT 94.935 93.190 95.105 93.360 ;
        RECT 94.935 92.830 95.105 93.000 ;
        RECT 94.935 92.470 95.105 92.640 ;
        RECT 88.545 92.110 88.715 92.280 ;
        RECT 89.340 92.150 89.510 92.320 ;
        RECT 93.710 92.150 93.880 92.320 ;
        RECT 94.070 92.150 94.240 92.320 ;
        RECT 88.545 91.750 88.715 91.920 ;
        RECT 94.935 92.110 95.105 92.280 ;
        RECT 88.545 91.390 88.715 91.560 ;
        RECT 88.545 91.030 88.715 91.200 ;
        RECT 88.545 90.670 88.715 90.840 ;
        RECT 88.545 90.310 88.715 90.480 ;
        RECT 89.925 91.730 90.095 91.900 ;
        RECT 89.925 91.370 90.095 91.540 ;
        RECT 89.925 91.010 90.095 91.180 ;
        RECT 89.925 90.650 90.095 90.820 ;
        RECT 89.925 90.290 90.095 90.460 ;
        RECT 93.055 91.730 93.225 91.900 ;
        RECT 93.055 91.370 93.225 91.540 ;
        RECT 93.055 91.010 93.225 91.180 ;
        RECT 93.055 90.650 93.225 90.820 ;
        RECT 93.055 90.290 93.225 90.460 ;
        RECT 94.935 91.750 95.105 91.920 ;
        RECT 94.935 91.390 95.105 91.560 ;
        RECT 94.935 91.030 95.105 91.200 ;
        RECT 94.935 90.670 95.105 90.840 ;
        RECT 94.935 90.310 95.105 90.480 ;
        RECT 88.545 89.950 88.715 90.120 ;
        RECT 89.340 89.870 89.510 90.040 ;
        RECT 93.710 89.870 93.880 90.040 ;
        RECT 94.070 89.870 94.240 90.040 ;
        RECT 94.935 89.950 95.105 90.120 ;
        RECT 88.545 89.590 88.715 89.760 ;
        RECT 94.935 89.590 95.105 89.760 ;
        RECT 88.845 89.200 89.015 89.370 ;
        RECT 89.205 89.200 89.375 89.370 ;
        RECT 89.565 89.200 89.735 89.370 ;
        RECT 89.925 89.200 90.095 89.370 ;
        RECT 90.285 89.200 90.455 89.370 ;
        RECT 90.645 89.200 90.815 89.370 ;
        RECT 92.115 89.200 92.285 89.370 ;
        RECT 92.475 89.200 92.645 89.370 ;
        RECT 92.835 89.200 93.005 89.370 ;
        RECT 93.195 89.200 93.365 89.370 ;
        RECT 93.555 89.200 93.725 89.370 ;
        RECT 93.915 89.200 94.085 89.370 ;
        RECT 94.275 89.200 94.445 89.370 ;
        RECT 94.635 89.200 94.805 89.370 ;
        RECT 108.635 111.940 108.805 112.110 ;
        RECT 110.555 113.500 110.725 113.670 ;
        RECT 110.555 113.140 110.725 113.310 ;
        RECT 110.555 112.780 110.725 112.950 ;
        RECT 110.555 112.420 110.725 112.590 ;
        RECT 110.555 112.060 110.725 112.230 ;
        RECT 111.925 113.500 112.095 113.670 ;
        RECT 111.925 113.140 112.095 113.310 ;
        RECT 111.925 112.780 112.095 112.950 ;
        RECT 111.925 112.420 112.095 112.590 ;
        RECT 111.925 112.060 112.095 112.230 ;
        RECT 113.845 113.550 114.015 113.720 ;
        RECT 118.195 114.260 118.365 114.430 ;
        RECT 119.400 114.280 119.570 114.450 ;
        RECT 119.760 114.280 119.930 114.450 ;
        RECT 120.415 114.280 120.585 114.450 ;
        RECT 120.965 114.160 121.135 114.330 ;
        RECT 119.400 113.850 119.570 114.020 ;
        RECT 119.760 113.850 119.930 114.020 ;
        RECT 113.845 113.190 114.015 113.360 ;
        RECT 113.845 112.830 114.015 113.000 ;
        RECT 113.845 112.470 114.015 112.640 ;
        RECT 113.845 112.110 114.015 112.280 ;
        RECT 108.635 111.580 108.805 111.750 ;
        RECT 109.690 111.640 109.860 111.810 ;
        RECT 110.050 111.640 110.220 111.810 ;
        RECT 111.060 111.640 111.230 111.810 ;
        RECT 111.420 111.640 111.590 111.810 ;
        RECT 112.430 111.640 112.600 111.810 ;
        RECT 112.790 111.640 112.960 111.810 ;
        RECT 113.845 111.750 114.015 111.920 ;
        RECT 113.845 111.390 114.015 111.560 ;
        RECT 108.635 111.220 108.805 111.390 ;
        RECT 108.635 110.860 108.805 111.030 ;
        RECT 108.635 110.500 108.805 110.670 ;
        RECT 108.635 110.140 108.805 110.310 ;
        RECT 108.635 109.780 108.805 109.950 ;
        RECT 110.555 111.220 110.725 111.390 ;
        RECT 110.555 110.860 110.725 111.030 ;
        RECT 110.555 110.500 110.725 110.670 ;
        RECT 110.555 110.140 110.725 110.310 ;
        RECT 110.555 109.780 110.725 109.950 ;
        RECT 111.925 111.220 112.095 111.390 ;
        RECT 111.925 110.860 112.095 111.030 ;
        RECT 111.925 110.500 112.095 110.670 ;
        RECT 111.925 110.140 112.095 110.310 ;
        RECT 111.925 109.780 112.095 109.950 ;
        RECT 113.845 111.030 114.015 111.200 ;
        RECT 113.845 110.670 114.015 110.840 ;
        RECT 113.845 110.310 114.015 110.480 ;
        RECT 113.845 109.950 114.015 110.120 ;
        RECT 108.635 109.420 108.805 109.590 ;
        RECT 113.845 109.590 114.015 109.760 ;
        RECT 114.925 113.465 115.095 113.635 ;
        RECT 115.535 113.525 115.705 113.695 ;
        RECT 115.895 113.525 116.065 113.695 ;
        RECT 116.255 113.525 116.425 113.695 ;
        RECT 116.615 113.525 116.785 113.695 ;
        RECT 116.975 113.525 117.145 113.695 ;
        RECT 117.335 113.525 117.505 113.695 ;
        RECT 114.925 113.105 115.095 113.275 ;
        RECT 114.925 112.745 115.095 112.915 ;
        RECT 115.980 112.855 116.150 113.025 ;
        RECT 116.340 112.855 116.510 113.025 ;
        RECT 117.395 112.905 117.565 113.075 ;
        RECT 114.925 112.385 115.095 112.555 ;
        RECT 115.475 112.425 115.645 112.595 ;
        RECT 115.980 112.425 116.150 112.595 ;
        RECT 116.340 112.425 116.510 112.595 ;
        RECT 117.395 112.545 117.565 112.715 ;
        RECT 114.925 112.025 115.095 112.195 ;
        RECT 117.395 112.185 117.565 112.355 ;
        RECT 115.980 111.995 116.150 112.165 ;
        RECT 116.340 111.995 116.510 112.165 ;
        RECT 117.395 111.825 117.565 111.995 ;
        RECT 115.980 111.565 116.150 111.735 ;
        RECT 116.340 111.565 116.510 111.735 ;
        RECT 116.845 111.565 117.015 111.735 ;
        RECT 114.925 111.385 115.095 111.555 ;
        RECT 117.395 111.465 117.565 111.635 ;
        RECT 114.925 111.025 115.095 111.195 ;
        RECT 115.980 111.135 116.150 111.305 ;
        RECT 116.340 111.135 116.510 111.305 ;
        RECT 117.395 111.105 117.565 111.275 ;
        RECT 114.925 110.665 115.095 110.835 ;
        RECT 115.475 110.705 115.645 110.875 ;
        RECT 115.980 110.705 116.150 110.875 ;
        RECT 116.340 110.705 116.510 110.875 ;
        RECT 117.395 110.745 117.565 110.915 ;
        RECT 114.925 110.305 115.095 110.475 ;
        RECT 115.980 110.275 116.150 110.445 ;
        RECT 116.340 110.275 116.510 110.445 ;
        RECT 117.395 110.385 117.565 110.555 ;
        RECT 117.395 110.025 117.565 110.195 ;
        RECT 114.985 109.605 115.155 109.775 ;
        RECT 115.345 109.605 115.515 109.775 ;
        RECT 115.705 109.605 115.875 109.775 ;
        RECT 116.065 109.605 116.235 109.775 ;
        RECT 116.425 109.605 116.595 109.775 ;
        RECT 116.785 109.605 116.955 109.775 ;
        RECT 117.395 109.665 117.565 109.835 ;
        RECT 118.195 113.670 118.365 113.840 ;
        RECT 120.965 113.800 121.135 113.970 ;
        RECT 118.195 113.310 118.365 113.480 ;
        RECT 119.400 113.420 119.570 113.590 ;
        RECT 119.760 113.420 119.930 113.590 ;
        RECT 120.415 113.420 120.585 113.590 ;
        RECT 120.965 113.440 121.135 113.610 ;
        RECT 118.195 112.950 118.365 113.120 ;
        RECT 119.400 112.990 119.570 113.160 ;
        RECT 119.760 112.990 119.930 113.160 ;
        RECT 120.965 113.080 121.135 113.250 ;
        RECT 118.195 112.590 118.365 112.760 ;
        RECT 118.745 112.560 118.915 112.730 ;
        RECT 119.400 112.560 119.570 112.730 ;
        RECT 119.760 112.560 119.930 112.730 ;
        RECT 120.965 112.720 121.135 112.890 ;
        RECT 118.195 112.230 118.365 112.400 ;
        RECT 120.965 112.360 121.135 112.530 ;
        RECT 119.400 112.130 119.570 112.300 ;
        RECT 119.760 112.130 119.930 112.300 ;
        RECT 118.195 111.870 118.365 112.040 ;
        RECT 120.965 112.000 121.135 112.170 ;
        RECT 118.745 111.700 118.915 111.870 ;
        RECT 119.400 111.700 119.570 111.870 ;
        RECT 119.760 111.700 119.930 111.870 ;
        RECT 118.195 111.510 118.365 111.680 ;
        RECT 120.965 111.640 121.135 111.810 ;
        RECT 118.195 111.150 118.365 111.320 ;
        RECT 119.400 111.270 119.570 111.440 ;
        RECT 119.760 111.270 119.930 111.440 ;
        RECT 120.965 111.280 121.135 111.450 ;
        RECT 118.195 110.790 118.365 110.960 ;
        RECT 118.745 110.840 118.915 111.010 ;
        RECT 119.400 110.840 119.570 111.010 ;
        RECT 119.760 110.840 119.930 111.010 ;
        RECT 120.965 110.920 121.135 111.090 ;
        RECT 118.195 110.430 118.365 110.600 ;
        RECT 119.400 110.410 119.570 110.580 ;
        RECT 119.760 110.410 119.930 110.580 ;
        RECT 120.965 110.560 121.135 110.730 ;
        RECT 120.965 110.200 121.135 110.370 ;
        RECT 118.255 109.780 118.425 109.950 ;
        RECT 118.615 109.780 118.785 109.950 ;
        RECT 118.975 109.780 119.145 109.950 ;
        RECT 119.335 109.780 119.505 109.950 ;
        RECT 119.695 109.780 119.865 109.950 ;
        RECT 120.055 109.780 120.225 109.950 ;
        RECT 120.415 109.780 120.585 109.950 ;
        RECT 120.965 109.840 121.135 110.010 ;
        RECT 121.840 118.060 122.010 118.230 ;
        RECT 121.840 117.700 122.010 117.870 ;
        RECT 121.840 117.340 122.010 117.510 ;
        RECT 121.840 116.980 122.010 117.150 ;
        RECT 121.840 116.620 122.010 116.790 ;
        RECT 122.390 118.060 122.560 118.230 ;
        RECT 122.390 117.700 122.560 117.870 ;
        RECT 122.390 117.340 122.560 117.510 ;
        RECT 122.390 116.980 122.560 117.150 ;
        RECT 122.390 116.620 122.560 116.790 ;
        RECT 123.760 118.060 123.930 118.230 ;
        RECT 123.760 117.700 123.930 117.870 ;
        RECT 123.760 117.340 123.930 117.510 ;
        RECT 123.760 116.980 123.930 117.150 ;
        RECT 123.760 116.620 123.930 116.790 ;
        RECT 125.130 118.060 125.300 118.230 ;
        RECT 125.130 117.700 125.300 117.870 ;
        RECT 125.130 117.340 125.300 117.510 ;
        RECT 125.130 116.980 125.300 117.150 ;
        RECT 125.130 116.620 125.300 116.790 ;
        RECT 125.680 117.910 125.850 118.080 ;
        RECT 125.680 117.550 125.850 117.720 ;
        RECT 125.680 117.190 125.850 117.360 ;
        RECT 125.680 116.830 125.850 117.000 ;
        RECT 121.840 116.260 122.010 116.430 ;
        RECT 125.680 116.470 125.850 116.640 ;
        RECT 122.895 116.200 123.065 116.370 ;
        RECT 123.255 116.200 123.425 116.370 ;
        RECT 124.265 116.200 124.435 116.370 ;
        RECT 124.625 116.200 124.795 116.370 ;
        RECT 121.840 115.900 122.010 116.070 ;
        RECT 125.680 116.110 125.850 116.280 ;
        RECT 121.840 115.540 122.010 115.710 ;
        RECT 121.840 115.180 122.010 115.350 ;
        RECT 121.840 114.820 122.010 114.990 ;
        RECT 121.840 114.460 122.010 114.630 ;
        RECT 122.390 115.780 122.560 115.950 ;
        RECT 122.390 115.420 122.560 115.590 ;
        RECT 122.390 115.060 122.560 115.230 ;
        RECT 122.390 114.700 122.560 114.870 ;
        RECT 122.390 114.340 122.560 114.510 ;
        RECT 123.760 115.780 123.930 115.950 ;
        RECT 123.760 115.420 123.930 115.590 ;
        RECT 123.760 115.060 123.930 115.230 ;
        RECT 123.760 114.700 123.930 114.870 ;
        RECT 123.760 114.340 123.930 114.510 ;
        RECT 125.130 115.780 125.300 115.950 ;
        RECT 125.130 115.420 125.300 115.590 ;
        RECT 125.130 115.060 125.300 115.230 ;
        RECT 125.130 114.700 125.300 114.870 ;
        RECT 125.130 114.340 125.300 114.510 ;
        RECT 125.680 115.750 125.850 115.920 ;
        RECT 125.680 115.390 125.850 115.560 ;
        RECT 125.680 115.030 125.850 115.200 ;
        RECT 125.680 114.670 125.850 114.840 ;
        RECT 121.840 114.100 122.010 114.270 ;
        RECT 125.680 114.310 125.850 114.480 ;
        RECT 122.895 113.920 123.065 114.090 ;
        RECT 123.255 113.920 123.425 114.090 ;
        RECT 124.265 113.920 124.435 114.090 ;
        RECT 124.625 113.920 124.795 114.090 ;
        RECT 125.680 113.950 125.850 114.120 ;
        RECT 121.840 113.740 122.010 113.910 ;
        RECT 121.840 113.380 122.010 113.550 ;
        RECT 121.840 113.020 122.010 113.190 ;
        RECT 121.840 112.660 122.010 112.830 ;
        RECT 121.840 112.300 122.010 112.470 ;
        RECT 121.840 111.940 122.010 112.110 ;
        RECT 122.390 113.500 122.560 113.670 ;
        RECT 122.390 113.140 122.560 113.310 ;
        RECT 122.390 112.780 122.560 112.950 ;
        RECT 122.390 112.420 122.560 112.590 ;
        RECT 122.390 112.060 122.560 112.230 ;
        RECT 123.760 113.500 123.930 113.670 ;
        RECT 123.760 113.140 123.930 113.310 ;
        RECT 123.760 112.780 123.930 112.950 ;
        RECT 123.760 112.420 123.930 112.590 ;
        RECT 123.760 112.060 123.930 112.230 ;
        RECT 125.130 113.500 125.300 113.670 ;
        RECT 125.130 113.140 125.300 113.310 ;
        RECT 125.130 112.780 125.300 112.950 ;
        RECT 125.130 112.420 125.300 112.590 ;
        RECT 125.130 112.060 125.300 112.230 ;
        RECT 125.680 113.590 125.850 113.760 ;
        RECT 125.680 113.230 125.850 113.400 ;
        RECT 125.680 112.870 125.850 113.040 ;
        RECT 125.680 112.510 125.850 112.680 ;
        RECT 125.680 112.150 125.850 112.320 ;
        RECT 121.840 111.580 122.010 111.750 ;
        RECT 122.895 111.640 123.065 111.810 ;
        RECT 123.255 111.640 123.425 111.810 ;
        RECT 124.265 111.640 124.435 111.810 ;
        RECT 124.625 111.640 124.795 111.810 ;
        RECT 125.680 111.790 125.850 111.960 ;
        RECT 125.680 111.430 125.850 111.600 ;
        RECT 121.840 111.220 122.010 111.390 ;
        RECT 121.840 110.860 122.010 111.030 ;
        RECT 121.840 110.500 122.010 110.670 ;
        RECT 121.840 110.140 122.010 110.310 ;
        RECT 121.840 109.780 122.010 109.950 ;
        RECT 122.390 111.220 122.560 111.390 ;
        RECT 122.390 110.860 122.560 111.030 ;
        RECT 122.390 110.500 122.560 110.670 ;
        RECT 122.390 110.140 122.560 110.310 ;
        RECT 122.390 109.780 122.560 109.950 ;
        RECT 123.760 111.220 123.930 111.390 ;
        RECT 123.760 110.860 123.930 111.030 ;
        RECT 123.760 110.500 123.930 110.670 ;
        RECT 123.760 110.140 123.930 110.310 ;
        RECT 123.760 109.780 123.930 109.950 ;
        RECT 125.130 111.220 125.300 111.390 ;
        RECT 125.130 110.860 125.300 111.030 ;
        RECT 125.130 110.500 125.300 110.670 ;
        RECT 125.130 110.140 125.300 110.310 ;
        RECT 125.130 109.780 125.300 109.950 ;
        RECT 125.680 111.070 125.850 111.240 ;
        RECT 125.680 110.710 125.850 110.880 ;
        RECT 125.680 110.350 125.850 110.520 ;
        RECT 125.680 109.990 125.850 110.160 ;
        RECT 109.690 109.360 109.860 109.530 ;
        RECT 110.050 109.360 110.220 109.530 ;
        RECT 111.060 109.360 111.230 109.530 ;
        RECT 111.420 109.360 111.590 109.530 ;
        RECT 112.430 109.360 112.600 109.530 ;
        RECT 112.790 109.360 112.960 109.530 ;
        RECT 108.635 109.060 108.805 109.230 ;
        RECT 113.845 109.230 114.015 109.400 ;
        RECT 108.635 108.700 108.805 108.870 ;
        RECT 108.635 108.340 108.805 108.510 ;
        RECT 108.635 107.980 108.805 108.150 ;
        RECT 108.635 107.620 108.805 107.790 ;
        RECT 110.555 108.940 110.725 109.110 ;
        RECT 110.555 108.580 110.725 108.750 ;
        RECT 110.555 108.220 110.725 108.390 ;
        RECT 110.555 107.860 110.725 108.030 ;
        RECT 110.555 107.500 110.725 107.670 ;
        RECT 111.925 108.940 112.095 109.110 ;
        RECT 111.925 108.580 112.095 108.750 ;
        RECT 111.925 108.220 112.095 108.390 ;
        RECT 111.925 107.860 112.095 108.030 ;
        RECT 111.925 107.500 112.095 107.670 ;
        RECT 113.845 108.870 114.015 109.040 ;
        RECT 113.845 108.510 114.015 108.680 ;
        RECT 113.845 108.150 114.015 108.320 ;
        RECT 113.845 107.790 114.015 107.960 ;
        RECT 108.635 107.260 108.805 107.430 ;
        RECT 113.845 107.430 114.015 107.600 ;
        RECT 109.690 107.080 109.860 107.250 ;
        RECT 110.050 107.080 110.220 107.250 ;
        RECT 111.060 107.080 111.230 107.250 ;
        RECT 111.420 107.080 111.590 107.250 ;
        RECT 112.430 107.080 112.600 107.250 ;
        RECT 112.790 107.080 112.960 107.250 ;
        RECT 108.635 106.900 108.805 107.070 ;
        RECT 113.845 107.070 114.015 107.240 ;
        RECT 108.635 106.540 108.805 106.710 ;
        RECT 108.635 106.180 108.805 106.350 ;
        RECT 108.635 105.820 108.805 105.990 ;
        RECT 108.635 105.460 108.805 105.630 ;
        RECT 108.635 105.100 108.805 105.270 ;
        RECT 110.555 106.660 110.725 106.830 ;
        RECT 110.555 106.300 110.725 106.470 ;
        RECT 110.555 105.940 110.725 106.110 ;
        RECT 110.555 105.580 110.725 105.750 ;
        RECT 110.555 105.220 110.725 105.390 ;
        RECT 111.925 106.660 112.095 106.830 ;
        RECT 111.925 106.300 112.095 106.470 ;
        RECT 111.925 105.940 112.095 106.110 ;
        RECT 111.925 105.580 112.095 105.750 ;
        RECT 111.925 105.220 112.095 105.390 ;
        RECT 113.845 106.710 114.015 106.880 ;
        RECT 113.845 106.350 114.015 106.520 ;
        RECT 113.845 105.990 114.015 106.160 ;
        RECT 113.845 105.630 114.015 105.800 ;
        RECT 113.845 105.270 114.015 105.440 ;
        RECT 108.635 104.740 108.805 104.910 ;
        RECT 109.690 104.800 109.860 104.970 ;
        RECT 110.050 104.800 110.220 104.970 ;
        RECT 111.060 104.800 111.230 104.970 ;
        RECT 111.420 104.800 111.590 104.970 ;
        RECT 112.430 104.800 112.600 104.970 ;
        RECT 112.790 104.800 112.960 104.970 ;
        RECT 113.845 104.910 114.015 105.080 ;
        RECT 113.845 104.550 114.015 104.720 ;
        RECT 108.635 104.380 108.805 104.550 ;
        RECT 108.635 104.020 108.805 104.190 ;
        RECT 108.635 103.660 108.805 103.830 ;
        RECT 108.635 103.300 108.805 103.470 ;
        RECT 108.635 102.940 108.805 103.110 ;
        RECT 110.555 104.380 110.725 104.550 ;
        RECT 110.555 104.020 110.725 104.190 ;
        RECT 110.555 103.660 110.725 103.830 ;
        RECT 110.555 103.300 110.725 103.470 ;
        RECT 110.555 102.940 110.725 103.110 ;
        RECT 111.925 104.380 112.095 104.550 ;
        RECT 111.925 104.020 112.095 104.190 ;
        RECT 111.925 103.660 112.095 103.830 ;
        RECT 111.925 103.300 112.095 103.470 ;
        RECT 111.925 102.940 112.095 103.110 ;
        RECT 113.845 104.190 114.015 104.360 ;
        RECT 113.845 103.830 114.015 104.000 ;
        RECT 113.845 103.470 114.015 103.640 ;
        RECT 113.845 103.110 114.015 103.280 ;
        RECT 108.635 102.580 108.805 102.750 ;
        RECT 113.845 102.750 114.015 102.920 ;
        RECT 109.690 102.520 109.860 102.690 ;
        RECT 110.050 102.520 110.220 102.690 ;
        RECT 111.060 102.520 111.230 102.690 ;
        RECT 111.420 102.520 111.590 102.690 ;
        RECT 112.430 102.520 112.600 102.690 ;
        RECT 112.790 102.520 112.960 102.690 ;
        RECT 108.635 102.220 108.805 102.390 ;
        RECT 113.845 102.390 114.015 102.560 ;
        RECT 108.635 101.860 108.805 102.030 ;
        RECT 108.635 101.500 108.805 101.670 ;
        RECT 108.635 101.140 108.805 101.310 ;
        RECT 108.635 100.780 108.805 100.950 ;
        RECT 110.555 102.100 110.725 102.270 ;
        RECT 110.555 101.740 110.725 101.910 ;
        RECT 110.555 101.380 110.725 101.550 ;
        RECT 110.555 101.020 110.725 101.190 ;
        RECT 110.555 100.660 110.725 100.830 ;
        RECT 111.925 102.100 112.095 102.270 ;
        RECT 111.925 101.740 112.095 101.910 ;
        RECT 111.925 101.380 112.095 101.550 ;
        RECT 111.925 101.020 112.095 101.190 ;
        RECT 111.925 100.660 112.095 100.830 ;
        RECT 113.845 102.030 114.015 102.200 ;
        RECT 113.845 101.670 114.015 101.840 ;
        RECT 113.845 101.310 114.015 101.480 ;
        RECT 113.845 100.950 114.015 101.120 ;
        RECT 108.635 100.420 108.805 100.590 ;
        RECT 113.845 100.590 114.015 100.760 ;
        RECT 109.690 100.240 109.860 100.410 ;
        RECT 110.050 100.240 110.220 100.410 ;
        RECT 111.060 100.240 111.230 100.410 ;
        RECT 111.420 100.240 111.590 100.410 ;
        RECT 112.430 100.240 112.600 100.410 ;
        RECT 112.790 100.240 112.960 100.410 ;
        RECT 108.635 100.060 108.805 100.230 ;
        RECT 113.845 100.230 114.015 100.400 ;
        RECT 108.635 99.700 108.805 99.870 ;
        RECT 108.635 99.340 108.805 99.510 ;
        RECT 108.635 98.980 108.805 99.150 ;
        RECT 108.635 98.620 108.805 98.790 ;
        RECT 108.635 98.260 108.805 98.430 ;
        RECT 110.555 99.820 110.725 99.990 ;
        RECT 110.555 99.460 110.725 99.630 ;
        RECT 110.555 99.100 110.725 99.270 ;
        RECT 110.555 98.740 110.725 98.910 ;
        RECT 110.555 98.380 110.725 98.550 ;
        RECT 111.925 99.820 112.095 99.990 ;
        RECT 111.925 99.460 112.095 99.630 ;
        RECT 111.925 99.100 112.095 99.270 ;
        RECT 111.925 98.740 112.095 98.910 ;
        RECT 111.925 98.380 112.095 98.550 ;
        RECT 113.845 99.870 114.015 100.040 ;
        RECT 113.845 99.510 114.015 99.680 ;
        RECT 113.845 99.150 114.015 99.320 ;
        RECT 113.845 98.790 114.015 98.960 ;
        RECT 113.845 98.430 114.015 98.600 ;
        RECT 108.635 97.900 108.805 98.070 ;
        RECT 109.690 97.960 109.860 98.130 ;
        RECT 110.050 97.960 110.220 98.130 ;
        RECT 111.060 97.960 111.230 98.130 ;
        RECT 111.420 97.960 111.590 98.130 ;
        RECT 112.430 97.960 112.600 98.130 ;
        RECT 112.790 97.960 112.960 98.130 ;
        RECT 113.845 98.070 114.015 98.240 ;
        RECT 113.845 97.710 114.015 97.880 ;
        RECT 108.635 97.540 108.805 97.710 ;
        RECT 108.635 97.180 108.805 97.350 ;
        RECT 108.635 96.820 108.805 96.990 ;
        RECT 108.635 96.460 108.805 96.630 ;
        RECT 108.635 96.100 108.805 96.270 ;
        RECT 110.555 97.540 110.725 97.710 ;
        RECT 110.555 97.180 110.725 97.350 ;
        RECT 110.555 96.820 110.725 96.990 ;
        RECT 110.555 96.460 110.725 96.630 ;
        RECT 110.555 96.100 110.725 96.270 ;
        RECT 111.925 97.540 112.095 97.710 ;
        RECT 111.925 97.180 112.095 97.350 ;
        RECT 111.925 96.820 112.095 96.990 ;
        RECT 111.925 96.460 112.095 96.630 ;
        RECT 111.925 96.100 112.095 96.270 ;
        RECT 113.845 97.350 114.015 97.520 ;
        RECT 113.845 96.990 114.015 97.160 ;
        RECT 113.845 96.630 114.015 96.800 ;
        RECT 113.845 96.270 114.015 96.440 ;
        RECT 108.635 95.740 108.805 95.910 ;
        RECT 113.845 95.910 114.015 96.080 ;
        RECT 109.690 95.680 109.860 95.850 ;
        RECT 110.050 95.680 110.220 95.850 ;
        RECT 111.060 95.680 111.230 95.850 ;
        RECT 111.420 95.680 111.590 95.850 ;
        RECT 112.430 95.680 112.600 95.850 ;
        RECT 112.790 95.680 112.960 95.850 ;
        RECT 108.635 95.380 108.805 95.550 ;
        RECT 113.845 95.550 114.015 95.720 ;
        RECT 108.635 95.020 108.805 95.190 ;
        RECT 108.635 94.660 108.805 94.830 ;
        RECT 108.635 94.300 108.805 94.470 ;
        RECT 108.635 93.940 108.805 94.110 ;
        RECT 110.555 95.260 110.725 95.430 ;
        RECT 110.555 94.900 110.725 95.070 ;
        RECT 110.555 94.540 110.725 94.710 ;
        RECT 110.555 94.180 110.725 94.350 ;
        RECT 110.555 93.820 110.725 93.990 ;
        RECT 111.925 95.260 112.095 95.430 ;
        RECT 111.925 94.900 112.095 95.070 ;
        RECT 111.925 94.540 112.095 94.710 ;
        RECT 111.925 94.180 112.095 94.350 ;
        RECT 111.925 93.820 112.095 93.990 ;
        RECT 113.845 95.190 114.015 95.360 ;
        RECT 113.845 94.830 114.015 95.000 ;
        RECT 113.845 94.470 114.015 94.640 ;
        RECT 113.845 94.110 114.015 94.280 ;
        RECT 108.635 93.580 108.805 93.750 ;
        RECT 113.845 93.750 114.015 93.920 ;
        RECT 109.690 93.400 109.860 93.570 ;
        RECT 110.050 93.400 110.220 93.570 ;
        RECT 111.060 93.400 111.230 93.570 ;
        RECT 111.420 93.400 111.590 93.570 ;
        RECT 112.430 93.400 112.600 93.570 ;
        RECT 112.790 93.400 112.960 93.570 ;
        RECT 108.635 93.220 108.805 93.390 ;
        RECT 113.845 93.390 114.015 93.560 ;
        RECT 108.635 92.860 108.805 93.030 ;
        RECT 108.635 92.500 108.805 92.670 ;
        RECT 108.635 92.140 108.805 92.310 ;
        RECT 108.635 91.780 108.805 91.950 ;
        RECT 108.635 91.420 108.805 91.590 ;
        RECT 110.555 92.980 110.725 93.150 ;
        RECT 110.555 92.620 110.725 92.790 ;
        RECT 110.555 92.260 110.725 92.430 ;
        RECT 110.555 91.900 110.725 92.070 ;
        RECT 110.555 91.540 110.725 91.710 ;
        RECT 111.925 92.980 112.095 93.150 ;
        RECT 111.925 92.620 112.095 92.790 ;
        RECT 111.925 92.260 112.095 92.430 ;
        RECT 111.925 91.900 112.095 92.070 ;
        RECT 111.925 91.540 112.095 91.710 ;
        RECT 113.845 93.030 114.015 93.200 ;
        RECT 113.845 92.670 114.015 92.840 ;
        RECT 113.845 92.310 114.015 92.480 ;
        RECT 113.845 91.950 114.015 92.120 ;
        RECT 113.845 91.590 114.015 91.760 ;
        RECT 108.635 91.060 108.805 91.230 ;
        RECT 109.690 91.120 109.860 91.290 ;
        RECT 110.050 91.120 110.220 91.290 ;
        RECT 111.060 91.120 111.230 91.290 ;
        RECT 111.420 91.120 111.590 91.290 ;
        RECT 112.430 91.120 112.600 91.290 ;
        RECT 112.790 91.120 112.960 91.290 ;
        RECT 113.845 91.230 114.015 91.400 ;
        RECT 113.845 90.870 114.015 91.040 ;
        RECT 108.635 90.700 108.805 90.870 ;
        RECT 108.635 90.340 108.805 90.510 ;
        RECT 108.635 89.980 108.805 90.150 ;
        RECT 108.635 89.620 108.805 89.790 ;
        RECT 108.635 89.260 108.805 89.430 ;
        RECT 110.555 90.700 110.725 90.870 ;
        RECT 110.555 90.340 110.725 90.510 ;
        RECT 110.555 89.980 110.725 90.150 ;
        RECT 110.555 89.620 110.725 89.790 ;
        RECT 110.555 89.260 110.725 89.430 ;
        RECT 111.925 90.700 112.095 90.870 ;
        RECT 111.925 90.340 112.095 90.510 ;
        RECT 111.925 89.980 112.095 90.150 ;
        RECT 111.925 89.620 112.095 89.790 ;
        RECT 111.925 89.260 112.095 89.430 ;
        RECT 113.845 90.510 114.015 90.680 ;
        RECT 113.845 90.150 114.015 90.320 ;
        RECT 113.845 89.790 114.015 89.960 ;
        RECT 113.845 89.430 114.015 89.600 ;
        RECT 108.635 88.900 108.805 89.070 ;
        RECT 113.845 89.070 114.015 89.240 ;
        RECT 109.690 88.840 109.860 89.010 ;
        RECT 110.050 88.840 110.220 89.010 ;
        RECT 111.060 88.840 111.230 89.010 ;
        RECT 111.420 88.840 111.590 89.010 ;
        RECT 112.430 88.840 112.600 89.010 ;
        RECT 112.790 88.840 112.960 89.010 ;
        RECT 108.635 88.540 108.805 88.710 ;
        RECT 113.845 88.710 114.015 88.880 ;
        RECT 108.635 88.180 108.805 88.350 ;
        RECT 108.635 87.820 108.805 87.990 ;
        RECT 108.635 87.460 108.805 87.630 ;
        RECT 108.635 87.100 108.805 87.270 ;
        RECT 110.555 88.420 110.725 88.590 ;
        RECT 110.555 88.060 110.725 88.230 ;
        RECT 110.555 87.700 110.725 87.870 ;
        RECT 110.555 87.340 110.725 87.510 ;
        RECT 110.555 86.980 110.725 87.150 ;
        RECT 111.925 88.420 112.095 88.590 ;
        RECT 111.925 88.060 112.095 88.230 ;
        RECT 111.925 87.700 112.095 87.870 ;
        RECT 111.925 87.340 112.095 87.510 ;
        RECT 111.925 86.980 112.095 87.150 ;
        RECT 113.845 88.350 114.015 88.520 ;
        RECT 113.845 87.990 114.015 88.160 ;
        RECT 113.845 87.630 114.015 87.800 ;
        RECT 113.845 87.270 114.015 87.440 ;
        RECT 108.635 86.740 108.805 86.910 ;
        RECT 113.845 86.910 114.015 87.080 ;
        RECT 109.690 86.560 109.860 86.730 ;
        RECT 110.050 86.560 110.220 86.730 ;
        RECT 111.060 86.560 111.230 86.730 ;
        RECT 111.420 86.560 111.590 86.730 ;
        RECT 112.430 86.560 112.600 86.730 ;
        RECT 112.790 86.560 112.960 86.730 ;
        RECT 108.635 86.380 108.805 86.550 ;
        RECT 113.845 86.550 114.015 86.720 ;
        RECT 108.635 86.020 108.805 86.190 ;
        RECT 108.635 85.660 108.805 85.830 ;
        RECT 108.635 85.300 108.805 85.470 ;
        RECT 108.635 84.940 108.805 85.110 ;
        RECT 108.635 84.580 108.805 84.750 ;
        RECT 110.555 86.140 110.725 86.310 ;
        RECT 110.555 85.780 110.725 85.950 ;
        RECT 110.555 85.420 110.725 85.590 ;
        RECT 110.555 85.060 110.725 85.230 ;
        RECT 110.555 84.700 110.725 84.870 ;
        RECT 111.925 86.140 112.095 86.310 ;
        RECT 111.925 85.780 112.095 85.950 ;
        RECT 111.925 85.420 112.095 85.590 ;
        RECT 111.925 85.060 112.095 85.230 ;
        RECT 111.925 84.700 112.095 84.870 ;
        RECT 113.845 86.190 114.015 86.360 ;
        RECT 113.845 85.830 114.015 86.000 ;
        RECT 113.845 85.470 114.015 85.640 ;
        RECT 113.845 85.110 114.015 85.280 ;
        RECT 113.845 84.750 114.015 84.920 ;
        RECT 108.635 84.220 108.805 84.390 ;
        RECT 109.690 84.280 109.860 84.450 ;
        RECT 110.050 84.280 110.220 84.450 ;
        RECT 111.060 84.280 111.230 84.450 ;
        RECT 111.420 84.280 111.590 84.450 ;
        RECT 112.430 84.280 112.600 84.450 ;
        RECT 112.790 84.280 112.960 84.450 ;
        RECT 113.845 84.390 114.015 84.560 ;
        RECT 113.845 84.030 114.015 84.200 ;
        RECT 121.840 109.420 122.010 109.590 ;
        RECT 125.680 109.630 125.850 109.800 ;
        RECT 122.895 109.360 123.065 109.530 ;
        RECT 123.255 109.360 123.425 109.530 ;
        RECT 124.265 109.360 124.435 109.530 ;
        RECT 124.625 109.360 124.795 109.530 ;
        RECT 121.840 109.060 122.010 109.230 ;
        RECT 125.680 109.270 125.850 109.440 ;
        RECT 121.840 108.700 122.010 108.870 ;
        RECT 121.840 108.340 122.010 108.510 ;
        RECT 121.840 107.980 122.010 108.150 ;
        RECT 121.840 107.620 122.010 107.790 ;
        RECT 122.390 108.940 122.560 109.110 ;
        RECT 122.390 108.580 122.560 108.750 ;
        RECT 122.390 108.220 122.560 108.390 ;
        RECT 122.390 107.860 122.560 108.030 ;
        RECT 122.390 107.500 122.560 107.670 ;
        RECT 123.760 108.940 123.930 109.110 ;
        RECT 123.760 108.580 123.930 108.750 ;
        RECT 123.760 108.220 123.930 108.390 ;
        RECT 123.760 107.860 123.930 108.030 ;
        RECT 123.760 107.500 123.930 107.670 ;
        RECT 125.130 108.940 125.300 109.110 ;
        RECT 125.130 108.580 125.300 108.750 ;
        RECT 125.130 108.220 125.300 108.390 ;
        RECT 125.130 107.860 125.300 108.030 ;
        RECT 125.130 107.500 125.300 107.670 ;
        RECT 125.680 108.910 125.850 109.080 ;
        RECT 125.680 108.550 125.850 108.720 ;
        RECT 125.680 108.190 125.850 108.360 ;
        RECT 125.680 107.830 125.850 108.000 ;
        RECT 121.840 107.260 122.010 107.430 ;
        RECT 125.680 107.470 125.850 107.640 ;
        RECT 122.895 107.080 123.065 107.250 ;
        RECT 123.255 107.080 123.425 107.250 ;
        RECT 124.265 107.080 124.435 107.250 ;
        RECT 124.625 107.080 124.795 107.250 ;
        RECT 125.680 107.110 125.850 107.280 ;
        RECT 121.840 106.900 122.010 107.070 ;
        RECT 121.840 106.540 122.010 106.710 ;
        RECT 121.840 106.180 122.010 106.350 ;
        RECT 121.840 105.820 122.010 105.990 ;
        RECT 121.840 105.460 122.010 105.630 ;
        RECT 121.840 105.100 122.010 105.270 ;
        RECT 122.390 106.660 122.560 106.830 ;
        RECT 122.390 106.300 122.560 106.470 ;
        RECT 122.390 105.940 122.560 106.110 ;
        RECT 122.390 105.580 122.560 105.750 ;
        RECT 122.390 105.220 122.560 105.390 ;
        RECT 123.760 106.660 123.930 106.830 ;
        RECT 123.760 106.300 123.930 106.470 ;
        RECT 123.760 105.940 123.930 106.110 ;
        RECT 123.760 105.580 123.930 105.750 ;
        RECT 123.760 105.220 123.930 105.390 ;
        RECT 125.130 106.660 125.300 106.830 ;
        RECT 125.130 106.300 125.300 106.470 ;
        RECT 125.130 105.940 125.300 106.110 ;
        RECT 125.130 105.580 125.300 105.750 ;
        RECT 125.130 105.220 125.300 105.390 ;
        RECT 125.680 106.750 125.850 106.920 ;
        RECT 125.680 106.390 125.850 106.560 ;
        RECT 125.680 106.030 125.850 106.200 ;
        RECT 125.680 105.670 125.850 105.840 ;
        RECT 125.680 105.310 125.850 105.480 ;
        RECT 121.840 104.740 122.010 104.910 ;
        RECT 122.895 104.800 123.065 104.970 ;
        RECT 123.255 104.800 123.425 104.970 ;
        RECT 124.265 104.800 124.435 104.970 ;
        RECT 124.625 104.800 124.795 104.970 ;
        RECT 125.680 104.950 125.850 105.120 ;
        RECT 125.680 104.590 125.850 104.760 ;
        RECT 121.840 104.380 122.010 104.550 ;
        RECT 121.840 104.020 122.010 104.190 ;
        RECT 121.840 103.660 122.010 103.830 ;
        RECT 121.840 103.300 122.010 103.470 ;
        RECT 121.840 102.940 122.010 103.110 ;
        RECT 122.390 104.380 122.560 104.550 ;
        RECT 122.390 104.020 122.560 104.190 ;
        RECT 122.390 103.660 122.560 103.830 ;
        RECT 122.390 103.300 122.560 103.470 ;
        RECT 122.390 102.940 122.560 103.110 ;
        RECT 123.760 104.380 123.930 104.550 ;
        RECT 123.760 104.020 123.930 104.190 ;
        RECT 123.760 103.660 123.930 103.830 ;
        RECT 123.760 103.300 123.930 103.470 ;
        RECT 123.760 102.940 123.930 103.110 ;
        RECT 125.130 104.380 125.300 104.550 ;
        RECT 125.130 104.020 125.300 104.190 ;
        RECT 125.130 103.660 125.300 103.830 ;
        RECT 125.130 103.300 125.300 103.470 ;
        RECT 125.130 102.940 125.300 103.110 ;
        RECT 125.680 104.230 125.850 104.400 ;
        RECT 125.680 103.870 125.850 104.040 ;
        RECT 125.680 103.510 125.850 103.680 ;
        RECT 125.680 103.150 125.850 103.320 ;
        RECT 121.840 102.580 122.010 102.750 ;
        RECT 125.680 102.790 125.850 102.960 ;
        RECT 122.895 102.520 123.065 102.690 ;
        RECT 123.255 102.520 123.425 102.690 ;
        RECT 124.265 102.520 124.435 102.690 ;
        RECT 124.625 102.520 124.795 102.690 ;
        RECT 121.840 102.220 122.010 102.390 ;
        RECT 125.680 102.430 125.850 102.600 ;
        RECT 121.840 101.860 122.010 102.030 ;
        RECT 121.840 101.500 122.010 101.670 ;
        RECT 121.840 101.140 122.010 101.310 ;
        RECT 121.840 100.780 122.010 100.950 ;
        RECT 122.390 102.100 122.560 102.270 ;
        RECT 122.390 101.740 122.560 101.910 ;
        RECT 122.390 101.380 122.560 101.550 ;
        RECT 122.390 101.020 122.560 101.190 ;
        RECT 122.390 100.660 122.560 100.830 ;
        RECT 123.760 102.100 123.930 102.270 ;
        RECT 123.760 101.740 123.930 101.910 ;
        RECT 123.760 101.380 123.930 101.550 ;
        RECT 123.760 101.020 123.930 101.190 ;
        RECT 123.760 100.660 123.930 100.830 ;
        RECT 125.130 102.100 125.300 102.270 ;
        RECT 125.130 101.740 125.300 101.910 ;
        RECT 125.130 101.380 125.300 101.550 ;
        RECT 125.130 101.020 125.300 101.190 ;
        RECT 125.130 100.660 125.300 100.830 ;
        RECT 125.680 102.070 125.850 102.240 ;
        RECT 125.680 101.710 125.850 101.880 ;
        RECT 125.680 101.350 125.850 101.520 ;
        RECT 125.680 100.990 125.850 101.160 ;
        RECT 121.840 100.420 122.010 100.590 ;
        RECT 125.680 100.630 125.850 100.800 ;
        RECT 122.895 100.240 123.065 100.410 ;
        RECT 123.255 100.240 123.425 100.410 ;
        RECT 124.265 100.240 124.435 100.410 ;
        RECT 124.625 100.240 124.795 100.410 ;
        RECT 125.680 100.270 125.850 100.440 ;
        RECT 121.840 100.060 122.010 100.230 ;
        RECT 121.840 99.700 122.010 99.870 ;
        RECT 121.840 99.340 122.010 99.510 ;
        RECT 121.840 98.980 122.010 99.150 ;
        RECT 121.840 98.620 122.010 98.790 ;
        RECT 121.840 98.260 122.010 98.430 ;
        RECT 122.390 99.820 122.560 99.990 ;
        RECT 122.390 99.460 122.560 99.630 ;
        RECT 122.390 99.100 122.560 99.270 ;
        RECT 122.390 98.740 122.560 98.910 ;
        RECT 122.390 98.380 122.560 98.550 ;
        RECT 123.760 99.820 123.930 99.990 ;
        RECT 123.760 99.460 123.930 99.630 ;
        RECT 123.760 99.100 123.930 99.270 ;
        RECT 123.760 98.740 123.930 98.910 ;
        RECT 123.760 98.380 123.930 98.550 ;
        RECT 125.130 99.820 125.300 99.990 ;
        RECT 125.130 99.460 125.300 99.630 ;
        RECT 125.130 99.100 125.300 99.270 ;
        RECT 125.130 98.740 125.300 98.910 ;
        RECT 125.130 98.380 125.300 98.550 ;
        RECT 125.680 99.910 125.850 100.080 ;
        RECT 125.680 99.550 125.850 99.720 ;
        RECT 125.680 99.190 125.850 99.360 ;
        RECT 125.680 98.830 125.850 99.000 ;
        RECT 125.680 98.470 125.850 98.640 ;
        RECT 121.840 97.900 122.010 98.070 ;
        RECT 122.895 97.960 123.065 98.130 ;
        RECT 123.255 97.960 123.425 98.130 ;
        RECT 124.265 97.960 124.435 98.130 ;
        RECT 124.625 97.960 124.795 98.130 ;
        RECT 125.680 98.110 125.850 98.280 ;
        RECT 125.680 97.750 125.850 97.920 ;
        RECT 121.840 97.540 122.010 97.710 ;
        RECT 121.840 97.180 122.010 97.350 ;
        RECT 121.840 96.820 122.010 96.990 ;
        RECT 121.840 96.460 122.010 96.630 ;
        RECT 121.840 96.100 122.010 96.270 ;
        RECT 122.390 97.540 122.560 97.710 ;
        RECT 122.390 97.180 122.560 97.350 ;
        RECT 122.390 96.820 122.560 96.990 ;
        RECT 122.390 96.460 122.560 96.630 ;
        RECT 122.390 96.100 122.560 96.270 ;
        RECT 123.760 97.540 123.930 97.710 ;
        RECT 123.760 97.180 123.930 97.350 ;
        RECT 123.760 96.820 123.930 96.990 ;
        RECT 123.760 96.460 123.930 96.630 ;
        RECT 123.760 96.100 123.930 96.270 ;
        RECT 125.130 97.540 125.300 97.710 ;
        RECT 125.130 97.180 125.300 97.350 ;
        RECT 125.130 96.820 125.300 96.990 ;
        RECT 125.130 96.460 125.300 96.630 ;
        RECT 125.130 96.100 125.300 96.270 ;
        RECT 125.680 97.390 125.850 97.560 ;
        RECT 125.680 97.030 125.850 97.200 ;
        RECT 125.680 96.670 125.850 96.840 ;
        RECT 125.680 96.310 125.850 96.480 ;
        RECT 121.840 95.740 122.010 95.910 ;
        RECT 125.680 95.950 125.850 96.120 ;
        RECT 122.895 95.680 123.065 95.850 ;
        RECT 123.255 95.680 123.425 95.850 ;
        RECT 124.265 95.680 124.435 95.850 ;
        RECT 124.625 95.680 124.795 95.850 ;
        RECT 121.840 95.380 122.010 95.550 ;
        RECT 125.680 95.590 125.850 95.760 ;
        RECT 121.840 95.020 122.010 95.190 ;
        RECT 121.840 94.660 122.010 94.830 ;
        RECT 121.840 94.300 122.010 94.470 ;
        RECT 121.840 93.940 122.010 94.110 ;
        RECT 122.390 95.260 122.560 95.430 ;
        RECT 122.390 94.900 122.560 95.070 ;
        RECT 122.390 94.540 122.560 94.710 ;
        RECT 122.390 94.180 122.560 94.350 ;
        RECT 122.390 93.820 122.560 93.990 ;
        RECT 123.760 95.260 123.930 95.430 ;
        RECT 123.760 94.900 123.930 95.070 ;
        RECT 123.760 94.540 123.930 94.710 ;
        RECT 123.760 94.180 123.930 94.350 ;
        RECT 123.760 93.820 123.930 93.990 ;
        RECT 125.130 95.260 125.300 95.430 ;
        RECT 125.130 94.900 125.300 95.070 ;
        RECT 125.130 94.540 125.300 94.710 ;
        RECT 125.130 94.180 125.300 94.350 ;
        RECT 125.130 93.820 125.300 93.990 ;
        RECT 125.680 95.230 125.850 95.400 ;
        RECT 125.680 94.870 125.850 95.040 ;
        RECT 125.680 94.510 125.850 94.680 ;
        RECT 125.680 94.150 125.850 94.320 ;
        RECT 121.840 93.580 122.010 93.750 ;
        RECT 125.680 93.790 125.850 93.960 ;
        RECT 122.895 93.400 123.065 93.570 ;
        RECT 123.255 93.400 123.425 93.570 ;
        RECT 124.265 93.400 124.435 93.570 ;
        RECT 124.625 93.400 124.795 93.570 ;
        RECT 125.680 93.430 125.850 93.600 ;
        RECT 121.840 93.220 122.010 93.390 ;
        RECT 121.840 92.860 122.010 93.030 ;
        RECT 121.840 92.500 122.010 92.670 ;
        RECT 121.840 92.140 122.010 92.310 ;
        RECT 121.840 91.780 122.010 91.950 ;
        RECT 121.840 91.420 122.010 91.590 ;
        RECT 122.390 92.980 122.560 93.150 ;
        RECT 122.390 92.620 122.560 92.790 ;
        RECT 122.390 92.260 122.560 92.430 ;
        RECT 122.390 91.900 122.560 92.070 ;
        RECT 122.390 91.540 122.560 91.710 ;
        RECT 123.760 92.980 123.930 93.150 ;
        RECT 123.760 92.620 123.930 92.790 ;
        RECT 123.760 92.260 123.930 92.430 ;
        RECT 123.760 91.900 123.930 92.070 ;
        RECT 123.760 91.540 123.930 91.710 ;
        RECT 125.130 92.980 125.300 93.150 ;
        RECT 125.130 92.620 125.300 92.790 ;
        RECT 125.130 92.260 125.300 92.430 ;
        RECT 125.130 91.900 125.300 92.070 ;
        RECT 125.130 91.540 125.300 91.710 ;
        RECT 125.680 93.070 125.850 93.240 ;
        RECT 125.680 92.710 125.850 92.880 ;
        RECT 125.680 92.350 125.850 92.520 ;
        RECT 125.680 91.990 125.850 92.160 ;
        RECT 125.680 91.630 125.850 91.800 ;
        RECT 121.840 91.060 122.010 91.230 ;
        RECT 122.895 91.120 123.065 91.290 ;
        RECT 123.255 91.120 123.425 91.290 ;
        RECT 124.265 91.120 124.435 91.290 ;
        RECT 124.625 91.120 124.795 91.290 ;
        RECT 125.680 91.270 125.850 91.440 ;
        RECT 125.680 90.910 125.850 91.080 ;
        RECT 121.840 90.700 122.010 90.870 ;
        RECT 121.840 90.340 122.010 90.510 ;
        RECT 121.840 89.980 122.010 90.150 ;
        RECT 121.840 89.620 122.010 89.790 ;
        RECT 121.840 89.260 122.010 89.430 ;
        RECT 122.390 90.700 122.560 90.870 ;
        RECT 122.390 90.340 122.560 90.510 ;
        RECT 122.390 89.980 122.560 90.150 ;
        RECT 122.390 89.620 122.560 89.790 ;
        RECT 122.390 89.260 122.560 89.430 ;
        RECT 125.130 90.700 125.300 90.870 ;
        RECT 125.130 90.340 125.300 90.510 ;
        RECT 125.130 89.980 125.300 90.150 ;
        RECT 125.130 89.620 125.300 89.790 ;
        RECT 125.130 89.260 125.300 89.430 ;
        RECT 125.680 90.550 125.850 90.720 ;
        RECT 125.680 90.190 125.850 90.360 ;
        RECT 125.680 89.830 125.850 90.000 ;
        RECT 125.680 89.470 125.850 89.640 ;
        RECT 121.840 88.900 122.010 89.070 ;
        RECT 125.680 89.110 125.850 89.280 ;
        RECT 122.895 88.840 123.065 89.010 ;
        RECT 123.255 88.840 123.425 89.010 ;
        RECT 124.265 88.840 124.435 89.010 ;
        RECT 124.625 88.840 124.795 89.010 ;
        RECT 121.840 88.540 122.010 88.710 ;
        RECT 125.680 88.750 125.850 88.920 ;
        RECT 121.840 88.180 122.010 88.350 ;
        RECT 121.840 87.820 122.010 87.990 ;
        RECT 121.840 87.460 122.010 87.630 ;
        RECT 121.840 87.100 122.010 87.270 ;
        RECT 122.390 88.420 122.560 88.590 ;
        RECT 122.390 88.060 122.560 88.230 ;
        RECT 122.390 87.700 122.560 87.870 ;
        RECT 122.390 87.340 122.560 87.510 ;
        RECT 122.390 86.980 122.560 87.150 ;
        RECT 125.130 88.420 125.300 88.590 ;
        RECT 125.130 88.060 125.300 88.230 ;
        RECT 125.130 87.700 125.300 87.870 ;
        RECT 125.130 87.340 125.300 87.510 ;
        RECT 125.130 86.980 125.300 87.150 ;
        RECT 125.680 88.390 125.850 88.560 ;
        RECT 125.680 88.030 125.850 88.200 ;
        RECT 125.680 87.670 125.850 87.840 ;
        RECT 125.680 87.310 125.850 87.480 ;
        RECT 121.840 86.740 122.010 86.910 ;
        RECT 125.680 86.950 125.850 87.120 ;
        RECT 122.895 86.560 123.065 86.730 ;
        RECT 123.255 86.560 123.425 86.730 ;
        RECT 124.265 86.560 124.435 86.730 ;
        RECT 124.625 86.560 124.795 86.730 ;
        RECT 125.680 86.590 125.850 86.760 ;
        RECT 121.840 86.380 122.010 86.550 ;
        RECT 121.840 86.020 122.010 86.190 ;
        RECT 121.840 85.660 122.010 85.830 ;
        RECT 121.840 85.300 122.010 85.470 ;
        RECT 121.840 84.940 122.010 85.110 ;
        RECT 121.840 84.580 122.010 84.750 ;
        RECT 122.390 86.140 122.560 86.310 ;
        RECT 122.390 85.780 122.560 85.950 ;
        RECT 122.390 85.420 122.560 85.590 ;
        RECT 122.390 85.060 122.560 85.230 ;
        RECT 122.390 84.700 122.560 84.870 ;
        RECT 125.130 86.140 125.300 86.310 ;
        RECT 125.130 85.780 125.300 85.950 ;
        RECT 125.130 85.420 125.300 85.590 ;
        RECT 125.130 85.060 125.300 85.230 ;
        RECT 125.130 84.700 125.300 84.870 ;
        RECT 125.680 86.230 125.850 86.400 ;
        RECT 125.680 85.870 125.850 86.040 ;
        RECT 125.680 85.510 125.850 85.680 ;
        RECT 125.680 85.150 125.850 85.320 ;
        RECT 125.680 84.790 125.850 84.960 ;
        RECT 121.840 84.220 122.010 84.390 ;
        RECT 122.895 84.280 123.065 84.450 ;
        RECT 123.255 84.280 123.425 84.450 ;
        RECT 124.265 84.280 124.435 84.450 ;
        RECT 124.625 84.280 124.795 84.450 ;
        RECT 125.680 84.430 125.850 84.600 ;
        RECT 108.635 83.860 108.805 84.030 ;
        RECT 108.635 83.500 108.805 83.670 ;
        RECT 88.805 83.020 88.975 83.190 ;
        RECT 89.165 83.020 89.335 83.190 ;
        RECT 89.525 83.020 89.695 83.190 ;
        RECT 89.885 83.020 90.055 83.190 ;
        RECT 90.245 83.020 90.415 83.190 ;
        RECT 90.605 83.020 90.775 83.190 ;
        RECT 92.100 83.020 92.270 83.190 ;
        RECT 92.460 83.020 92.630 83.190 ;
        RECT 92.820 83.020 92.990 83.190 ;
        RECT 93.180 83.020 93.350 83.190 ;
        RECT 93.540 83.020 93.710 83.190 ;
        RECT 93.900 83.020 94.070 83.190 ;
        RECT 94.260 83.020 94.430 83.190 ;
        RECT 94.620 83.020 94.790 83.190 ;
        RECT 71.775 82.670 71.945 82.840 ;
        RECT 72.135 82.670 72.305 82.840 ;
        RECT 72.495 82.670 72.665 82.840 ;
        RECT 72.855 82.670 73.025 82.840 ;
        RECT 73.215 82.670 73.385 82.840 ;
        RECT 73.575 82.670 73.745 82.840 ;
        RECT 75.295 82.670 75.465 82.840 ;
        RECT 75.655 82.670 75.825 82.840 ;
        RECT 76.015 82.670 76.185 82.840 ;
        RECT 76.375 82.670 76.545 82.840 ;
        RECT 76.735 82.670 76.905 82.840 ;
        RECT 77.095 82.670 77.265 82.840 ;
        RECT 77.455 82.670 77.625 82.840 ;
        RECT 77.815 82.670 77.985 82.840 ;
        RECT 78.175 82.670 78.345 82.840 ;
        RECT 78.535 82.670 78.705 82.840 ;
        RECT 78.895 82.670 79.065 82.840 ;
        RECT 79.495 82.670 79.665 82.840 ;
        RECT 79.855 82.670 80.025 82.840 ;
        RECT 80.215 82.670 80.385 82.840 ;
        RECT 80.575 82.670 80.745 82.840 ;
        RECT 80.935 82.670 81.105 82.840 ;
        RECT 81.295 82.670 81.465 82.840 ;
        RECT 81.655 82.670 81.825 82.840 ;
        RECT 82.015 82.670 82.185 82.840 ;
        RECT 82.375 82.670 82.545 82.840 ;
        RECT 82.735 82.670 82.905 82.840 ;
        RECT 83.095 82.670 83.265 82.840 ;
        RECT 84.815 82.670 84.985 82.840 ;
        RECT 85.175 82.670 85.345 82.840 ;
        RECT 85.535 82.670 85.705 82.840 ;
        RECT 85.895 82.670 86.065 82.840 ;
        RECT 86.255 82.670 86.425 82.840 ;
        RECT 86.615 82.670 86.785 82.840 ;
        RECT 71.475 82.320 71.645 82.490 ;
        RECT 79.195 82.320 79.365 82.490 ;
        RECT 71.475 81.960 71.645 82.130 ;
        RECT 72.680 82.000 72.850 82.170 ;
        RECT 73.040 82.000 73.210 82.170 ;
        RECT 75.980 82.000 76.150 82.170 ;
        RECT 76.340 82.000 76.510 82.170 ;
        RECT 77.630 82.000 77.800 82.170 ;
        RECT 77.990 82.000 78.160 82.170 ;
        RECT 86.915 82.320 87.085 82.490 ;
        RECT 79.195 81.960 79.365 82.130 ;
        RECT 80.400 82.000 80.570 82.170 ;
        RECT 80.760 82.000 80.930 82.170 ;
        RECT 82.050 82.000 82.220 82.170 ;
        RECT 82.410 82.000 82.580 82.170 ;
        RECT 85.350 82.000 85.520 82.170 ;
        RECT 85.710 82.000 85.880 82.170 ;
        RECT 71.475 81.600 71.645 81.770 ;
        RECT 71.475 81.240 71.645 81.410 ;
        RECT 72.025 81.750 72.195 81.920 ;
        RECT 73.695 81.750 73.865 81.920 ;
        RECT 72.680 81.570 72.850 81.740 ;
        RECT 73.040 81.570 73.210 81.740 ;
        RECT 72.025 81.390 72.195 81.560 ;
        RECT 73.695 81.390 73.865 81.560 ;
        RECT 75.325 81.750 75.495 81.920 ;
        RECT 78.645 81.750 78.815 81.920 ;
        RECT 75.980 81.570 76.150 81.740 ;
        RECT 76.340 81.570 76.510 81.740 ;
        RECT 77.630 81.570 77.800 81.740 ;
        RECT 77.990 81.570 78.160 81.740 ;
        RECT 75.325 81.390 75.495 81.560 ;
        RECT 78.645 81.390 78.815 81.560 ;
        RECT 86.915 81.960 87.085 82.130 ;
        RECT 79.195 81.600 79.365 81.770 ;
        RECT 72.680 81.140 72.850 81.310 ;
        RECT 73.040 81.140 73.210 81.310 ;
        RECT 75.980 81.140 76.150 81.310 ;
        RECT 76.340 81.140 76.510 81.310 ;
        RECT 77.630 81.140 77.800 81.310 ;
        RECT 77.990 81.140 78.160 81.310 ;
        RECT 79.195 81.240 79.365 81.410 ;
        RECT 79.745 81.750 79.915 81.920 ;
        RECT 83.065 81.750 83.235 81.920 ;
        RECT 80.400 81.570 80.570 81.740 ;
        RECT 80.760 81.570 80.930 81.740 ;
        RECT 82.050 81.570 82.220 81.740 ;
        RECT 82.410 81.570 82.580 81.740 ;
        RECT 79.745 81.390 79.915 81.560 ;
        RECT 83.065 81.390 83.235 81.560 ;
        RECT 84.695 81.750 84.865 81.920 ;
        RECT 86.365 81.750 86.535 81.920 ;
        RECT 85.350 81.570 85.520 81.740 ;
        RECT 85.710 81.570 85.880 81.740 ;
        RECT 84.695 81.390 84.865 81.560 ;
        RECT 86.365 81.390 86.535 81.560 ;
        RECT 86.915 81.600 87.085 81.770 ;
        RECT 71.475 80.880 71.645 81.050 ;
        RECT 71.475 80.520 71.645 80.690 ;
        RECT 72.025 80.890 72.195 81.060 ;
        RECT 73.695 80.890 73.865 81.060 ;
        RECT 72.680 80.710 72.850 80.880 ;
        RECT 73.040 80.710 73.210 80.880 ;
        RECT 72.025 80.530 72.195 80.700 ;
        RECT 73.695 80.530 73.865 80.700 ;
        RECT 75.325 80.890 75.495 81.060 ;
        RECT 78.645 80.890 78.815 81.060 ;
        RECT 75.980 80.710 76.150 80.880 ;
        RECT 76.340 80.710 76.510 80.880 ;
        RECT 77.630 80.710 77.800 80.880 ;
        RECT 77.990 80.710 78.160 80.880 ;
        RECT 75.325 80.530 75.495 80.700 ;
        RECT 78.645 80.530 78.815 80.700 ;
        RECT 80.400 81.140 80.570 81.310 ;
        RECT 80.760 81.140 80.930 81.310 ;
        RECT 82.050 81.140 82.220 81.310 ;
        RECT 82.410 81.140 82.580 81.310 ;
        RECT 85.350 81.140 85.520 81.310 ;
        RECT 85.710 81.140 85.880 81.310 ;
        RECT 86.915 81.240 87.085 81.410 ;
        RECT 79.195 80.880 79.365 81.050 ;
        RECT 79.195 80.520 79.365 80.690 ;
        RECT 79.745 80.890 79.915 81.060 ;
        RECT 83.065 80.890 83.235 81.060 ;
        RECT 80.400 80.710 80.570 80.880 ;
        RECT 80.760 80.710 80.930 80.880 ;
        RECT 82.050 80.710 82.220 80.880 ;
        RECT 82.410 80.710 82.580 80.880 ;
        RECT 79.745 80.530 79.915 80.700 ;
        RECT 83.065 80.530 83.235 80.700 ;
        RECT 84.695 80.890 84.865 81.060 ;
        RECT 86.365 80.890 86.535 81.060 ;
        RECT 85.350 80.710 85.520 80.880 ;
        RECT 85.710 80.710 85.880 80.880 ;
        RECT 84.695 80.530 84.865 80.700 ;
        RECT 86.365 80.530 86.535 80.700 ;
        RECT 86.915 80.880 87.085 81.050 ;
        RECT 71.475 80.160 71.645 80.330 ;
        RECT 72.680 80.280 72.850 80.450 ;
        RECT 73.040 80.280 73.210 80.450 ;
        RECT 75.980 80.280 76.150 80.450 ;
        RECT 76.340 80.280 76.510 80.450 ;
        RECT 77.630 80.280 77.800 80.450 ;
        RECT 77.990 80.280 78.160 80.450 ;
        RECT 86.915 80.520 87.085 80.690 ;
        RECT 71.475 79.800 71.645 79.970 ;
        RECT 72.025 80.030 72.195 80.200 ;
        RECT 73.695 80.030 73.865 80.200 ;
        RECT 72.680 79.850 72.850 80.020 ;
        RECT 73.040 79.850 73.210 80.020 ;
        RECT 72.025 79.670 72.195 79.840 ;
        RECT 73.695 79.670 73.865 79.840 ;
        RECT 75.325 80.030 75.495 80.200 ;
        RECT 78.645 80.030 78.815 80.200 ;
        RECT 75.980 79.850 76.150 80.020 ;
        RECT 76.340 79.850 76.510 80.020 ;
        RECT 77.630 79.850 77.800 80.020 ;
        RECT 77.990 79.850 78.160 80.020 ;
        RECT 75.325 79.670 75.495 79.840 ;
        RECT 78.645 79.670 78.815 79.840 ;
        RECT 79.195 80.160 79.365 80.330 ;
        RECT 80.400 80.280 80.570 80.450 ;
        RECT 80.760 80.280 80.930 80.450 ;
        RECT 82.050 80.280 82.220 80.450 ;
        RECT 82.410 80.280 82.580 80.450 ;
        RECT 85.350 80.280 85.520 80.450 ;
        RECT 85.710 80.280 85.880 80.450 ;
        RECT 79.195 79.800 79.365 79.970 ;
        RECT 71.475 79.440 71.645 79.610 ;
        RECT 79.745 80.030 79.915 80.200 ;
        RECT 83.065 80.030 83.235 80.200 ;
        RECT 80.400 79.850 80.570 80.020 ;
        RECT 80.760 79.850 80.930 80.020 ;
        RECT 82.050 79.850 82.220 80.020 ;
        RECT 82.410 79.850 82.580 80.020 ;
        RECT 79.745 79.670 79.915 79.840 ;
        RECT 83.065 79.670 83.235 79.840 ;
        RECT 84.695 80.030 84.865 80.200 ;
        RECT 86.365 80.030 86.535 80.200 ;
        RECT 85.350 79.850 85.520 80.020 ;
        RECT 85.710 79.850 85.880 80.020 ;
        RECT 84.695 79.670 84.865 79.840 ;
        RECT 86.365 79.670 86.535 79.840 ;
        RECT 86.915 80.160 87.085 80.330 ;
        RECT 86.915 79.800 87.085 79.970 ;
        RECT 72.680 79.420 72.850 79.590 ;
        RECT 73.040 79.420 73.210 79.590 ;
        RECT 75.980 79.420 76.150 79.590 ;
        RECT 76.340 79.420 76.510 79.590 ;
        RECT 77.630 79.420 77.800 79.590 ;
        RECT 77.990 79.420 78.160 79.590 ;
        RECT 79.195 79.440 79.365 79.610 ;
        RECT 71.475 79.080 71.645 79.250 ;
        RECT 71.475 78.720 71.645 78.890 ;
        RECT 72.025 79.170 72.195 79.340 ;
        RECT 73.695 79.170 73.865 79.340 ;
        RECT 72.680 78.990 72.850 79.160 ;
        RECT 73.040 78.990 73.210 79.160 ;
        RECT 72.025 78.810 72.195 78.980 ;
        RECT 73.695 78.810 73.865 78.980 ;
        RECT 75.325 79.170 75.495 79.340 ;
        RECT 78.645 79.170 78.815 79.340 ;
        RECT 75.980 78.990 76.150 79.160 ;
        RECT 76.340 78.990 76.510 79.160 ;
        RECT 77.630 78.990 77.800 79.160 ;
        RECT 77.990 78.990 78.160 79.160 ;
        RECT 75.325 78.810 75.495 78.980 ;
        RECT 78.645 78.810 78.815 78.980 ;
        RECT 80.400 79.420 80.570 79.590 ;
        RECT 80.760 79.420 80.930 79.590 ;
        RECT 82.050 79.420 82.220 79.590 ;
        RECT 82.410 79.420 82.580 79.590 ;
        RECT 85.350 79.420 85.520 79.590 ;
        RECT 85.710 79.420 85.880 79.590 ;
        RECT 86.915 79.440 87.085 79.610 ;
        RECT 79.195 79.080 79.365 79.250 ;
        RECT 72.680 78.560 72.850 78.730 ;
        RECT 73.040 78.560 73.210 78.730 ;
        RECT 75.980 78.560 76.150 78.730 ;
        RECT 76.340 78.560 76.510 78.730 ;
        RECT 77.630 78.560 77.800 78.730 ;
        RECT 77.990 78.560 78.160 78.730 ;
        RECT 79.195 78.720 79.365 78.890 ;
        RECT 79.745 79.170 79.915 79.340 ;
        RECT 83.065 79.170 83.235 79.340 ;
        RECT 80.400 78.990 80.570 79.160 ;
        RECT 80.760 78.990 80.930 79.160 ;
        RECT 82.050 78.990 82.220 79.160 ;
        RECT 82.410 78.990 82.580 79.160 ;
        RECT 79.745 78.810 79.915 78.980 ;
        RECT 83.065 78.810 83.235 78.980 ;
        RECT 84.695 79.170 84.865 79.340 ;
        RECT 86.365 79.170 86.535 79.340 ;
        RECT 85.350 78.990 85.520 79.160 ;
        RECT 85.710 78.990 85.880 79.160 ;
        RECT 84.695 78.810 84.865 78.980 ;
        RECT 86.365 78.810 86.535 78.980 ;
        RECT 86.915 79.080 87.085 79.250 ;
        RECT 71.475 78.360 71.645 78.530 ;
        RECT 80.400 78.560 80.570 78.730 ;
        RECT 80.760 78.560 80.930 78.730 ;
        RECT 82.050 78.560 82.220 78.730 ;
        RECT 82.410 78.560 82.580 78.730 ;
        RECT 85.350 78.560 85.520 78.730 ;
        RECT 85.710 78.560 85.880 78.730 ;
        RECT 86.915 78.720 87.085 78.890 ;
        RECT 79.195 78.360 79.365 78.530 ;
        RECT 86.915 78.360 87.085 78.530 ;
        RECT 88.505 82.670 88.675 82.840 ;
        RECT 94.920 82.670 95.090 82.840 ;
        RECT 88.505 82.310 88.675 82.480 ;
        RECT 89.345 82.350 89.515 82.520 ;
        RECT 89.705 82.350 89.875 82.520 ;
        RECT 92.655 82.350 92.825 82.520 ;
        RECT 93.015 82.350 93.185 82.520 ;
        RECT 93.375 82.350 93.545 82.520 ;
        RECT 93.735 82.350 93.905 82.520 ;
        RECT 94.095 82.350 94.265 82.520 ;
        RECT 94.920 82.310 95.090 82.480 ;
        RECT 88.505 81.950 88.675 82.120 ;
        RECT 90.360 82.100 90.530 82.270 ;
        RECT 89.345 81.920 89.515 82.090 ;
        RECT 89.705 81.920 89.875 82.090 ;
        RECT 88.505 81.590 88.675 81.760 ;
        RECT 90.360 81.740 90.530 81.910 ;
        RECT 92.040 82.100 92.210 82.270 ;
        RECT 92.655 81.920 92.825 82.090 ;
        RECT 93.015 81.920 93.185 82.090 ;
        RECT 93.375 81.920 93.545 82.090 ;
        RECT 93.735 81.920 93.905 82.090 ;
        RECT 94.095 81.920 94.265 82.090 ;
        RECT 94.920 81.950 95.090 82.120 ;
        RECT 92.040 81.740 92.210 81.910 ;
        RECT 89.345 81.490 89.515 81.660 ;
        RECT 89.705 81.490 89.875 81.660 ;
        RECT 92.655 81.490 92.825 81.660 ;
        RECT 93.015 81.490 93.185 81.660 ;
        RECT 93.375 81.490 93.545 81.660 ;
        RECT 93.735 81.490 93.905 81.660 ;
        RECT 94.095 81.490 94.265 81.660 ;
        RECT 94.920 81.590 95.090 81.760 ;
        RECT 88.505 81.230 88.675 81.400 ;
        RECT 90.360 81.240 90.530 81.410 ;
        RECT 89.345 81.060 89.515 81.230 ;
        RECT 89.705 81.060 89.875 81.230 ;
        RECT 88.505 80.870 88.675 81.040 ;
        RECT 90.360 80.880 90.530 81.050 ;
        RECT 92.040 81.240 92.210 81.410 ;
        RECT 94.920 81.230 95.090 81.400 ;
        RECT 92.655 81.060 92.825 81.230 ;
        RECT 93.015 81.060 93.185 81.230 ;
        RECT 93.375 81.060 93.545 81.230 ;
        RECT 93.735 81.060 93.905 81.230 ;
        RECT 94.095 81.060 94.265 81.230 ;
        RECT 92.040 80.880 92.210 81.050 ;
        RECT 94.920 80.870 95.090 81.040 ;
        RECT 88.505 80.510 88.675 80.680 ;
        RECT 89.345 80.630 89.515 80.800 ;
        RECT 89.705 80.630 89.875 80.800 ;
        RECT 92.655 80.630 92.825 80.800 ;
        RECT 93.015 80.630 93.185 80.800 ;
        RECT 93.375 80.630 93.545 80.800 ;
        RECT 93.735 80.630 93.905 80.800 ;
        RECT 94.095 80.630 94.265 80.800 ;
        RECT 90.360 80.380 90.530 80.550 ;
        RECT 88.505 80.150 88.675 80.320 ;
        RECT 89.345 80.200 89.515 80.370 ;
        RECT 89.705 80.200 89.875 80.370 ;
        RECT 90.360 80.020 90.530 80.190 ;
        RECT 92.040 80.380 92.210 80.550 ;
        RECT 94.920 80.510 95.090 80.680 ;
        RECT 92.655 80.200 92.825 80.370 ;
        RECT 93.015 80.200 93.185 80.370 ;
        RECT 93.375 80.200 93.545 80.370 ;
        RECT 93.735 80.200 93.905 80.370 ;
        RECT 94.095 80.200 94.265 80.370 ;
        RECT 92.040 80.020 92.210 80.190 ;
        RECT 94.920 80.150 95.090 80.320 ;
        RECT 88.505 79.790 88.675 79.960 ;
        RECT 89.345 79.770 89.515 79.940 ;
        RECT 89.705 79.770 89.875 79.940 ;
        RECT 92.655 79.770 92.825 79.940 ;
        RECT 93.015 79.770 93.185 79.940 ;
        RECT 93.375 79.770 93.545 79.940 ;
        RECT 93.735 79.770 93.905 79.940 ;
        RECT 94.095 79.770 94.265 79.940 ;
        RECT 94.920 79.790 95.090 79.960 ;
        RECT 88.505 79.430 88.675 79.600 ;
        RECT 90.360 79.520 90.530 79.690 ;
        RECT 89.345 79.340 89.515 79.510 ;
        RECT 89.705 79.340 89.875 79.510 ;
        RECT 88.505 79.070 88.675 79.240 ;
        RECT 90.360 79.160 90.530 79.330 ;
        RECT 92.040 79.520 92.210 79.690 ;
        RECT 92.655 79.340 92.825 79.510 ;
        RECT 93.015 79.340 93.185 79.510 ;
        RECT 93.375 79.340 93.545 79.510 ;
        RECT 93.735 79.340 93.905 79.510 ;
        RECT 94.095 79.340 94.265 79.510 ;
        RECT 94.920 79.430 95.090 79.600 ;
        RECT 92.040 79.160 92.210 79.330 ;
        RECT 89.345 78.910 89.515 79.080 ;
        RECT 89.705 78.910 89.875 79.080 ;
        RECT 92.655 78.910 92.825 79.080 ;
        RECT 93.015 78.910 93.185 79.080 ;
        RECT 93.375 78.910 93.545 79.080 ;
        RECT 93.735 78.910 93.905 79.080 ;
        RECT 94.095 78.910 94.265 79.080 ;
        RECT 94.920 79.070 95.090 79.240 ;
        RECT 88.505 78.710 88.675 78.880 ;
        RECT 94.920 78.710 95.090 78.880 ;
        RECT 88.805 78.240 88.975 78.410 ;
        RECT 89.165 78.240 89.335 78.410 ;
        RECT 89.525 78.240 89.695 78.410 ;
        RECT 89.885 78.240 90.055 78.410 ;
        RECT 90.245 78.240 90.415 78.410 ;
        RECT 90.605 78.240 90.775 78.410 ;
        RECT 92.100 78.240 92.270 78.410 ;
        RECT 92.460 78.240 92.630 78.410 ;
        RECT 92.820 78.240 92.990 78.410 ;
        RECT 93.180 78.240 93.350 78.410 ;
        RECT 93.540 78.240 93.710 78.410 ;
        RECT 93.900 78.240 94.070 78.410 ;
        RECT 94.260 78.240 94.430 78.410 ;
        RECT 94.620 78.240 94.790 78.410 ;
        RECT 108.635 83.140 108.805 83.310 ;
        RECT 108.635 82.780 108.805 82.950 ;
        RECT 108.635 82.420 108.805 82.590 ;
        RECT 110.555 83.860 110.725 84.030 ;
        RECT 110.555 83.500 110.725 83.670 ;
        RECT 110.555 83.140 110.725 83.310 ;
        RECT 110.555 82.780 110.725 82.950 ;
        RECT 110.555 82.420 110.725 82.590 ;
        RECT 111.925 83.860 112.095 84.030 ;
        RECT 111.925 83.500 112.095 83.670 ;
        RECT 111.925 83.140 112.095 83.310 ;
        RECT 111.925 82.780 112.095 82.950 ;
        RECT 111.925 82.420 112.095 82.590 ;
        RECT 113.845 83.670 114.015 83.840 ;
        RECT 113.845 83.310 114.015 83.480 ;
        RECT 113.845 82.950 114.015 83.120 ;
        RECT 113.845 82.590 114.015 82.760 ;
        RECT 108.635 82.060 108.805 82.230 ;
        RECT 113.845 82.230 114.015 82.400 ;
        RECT 109.690 82.000 109.860 82.170 ;
        RECT 110.050 82.000 110.220 82.170 ;
        RECT 111.060 82.000 111.230 82.170 ;
        RECT 111.420 82.000 111.590 82.170 ;
        RECT 112.430 82.000 112.600 82.170 ;
        RECT 112.790 82.000 112.960 82.170 ;
        RECT 108.635 81.700 108.805 81.870 ;
        RECT 113.845 81.870 114.015 82.040 ;
        RECT 108.635 81.340 108.805 81.510 ;
        RECT 108.635 80.980 108.805 81.150 ;
        RECT 108.635 80.620 108.805 80.790 ;
        RECT 108.635 80.260 108.805 80.430 ;
        RECT 110.555 81.580 110.725 81.750 ;
        RECT 110.555 81.220 110.725 81.390 ;
        RECT 110.555 80.860 110.725 81.030 ;
        RECT 110.555 80.500 110.725 80.670 ;
        RECT 110.555 80.140 110.725 80.310 ;
        RECT 111.925 81.580 112.095 81.750 ;
        RECT 111.925 81.220 112.095 81.390 ;
        RECT 111.925 80.860 112.095 81.030 ;
        RECT 111.925 80.500 112.095 80.670 ;
        RECT 111.925 80.140 112.095 80.310 ;
        RECT 113.845 81.510 114.015 81.680 ;
        RECT 113.845 81.150 114.015 81.320 ;
        RECT 113.845 80.790 114.015 80.960 ;
        RECT 113.845 80.430 114.015 80.600 ;
        RECT 108.635 79.900 108.805 80.070 ;
        RECT 113.845 80.070 114.015 80.240 ;
        RECT 114.925 83.895 115.095 84.065 ;
        RECT 115.535 83.955 115.705 84.125 ;
        RECT 115.895 83.955 116.065 84.125 ;
        RECT 116.255 83.955 116.425 84.125 ;
        RECT 116.615 83.955 116.785 84.125 ;
        RECT 116.975 83.955 117.145 84.125 ;
        RECT 117.335 83.955 117.505 84.125 ;
        RECT 114.925 83.535 115.095 83.705 ;
        RECT 125.680 84.070 125.850 84.240 ;
        RECT 114.925 83.175 115.095 83.345 ;
        RECT 115.980 83.325 116.150 83.495 ;
        RECT 116.340 83.325 116.510 83.495 ;
        RECT 117.395 83.415 117.565 83.585 ;
        RECT 114.925 82.815 115.095 82.985 ;
        RECT 115.980 82.895 116.150 83.065 ;
        RECT 116.340 82.895 116.510 83.065 ;
        RECT 116.845 82.895 117.015 83.065 ;
        RECT 117.395 83.055 117.565 83.225 ;
        RECT 117.395 82.695 117.565 82.865 ;
        RECT 114.925 82.455 115.095 82.625 ;
        RECT 115.980 82.465 116.150 82.635 ;
        RECT 116.340 82.465 116.510 82.635 ;
        RECT 117.395 82.335 117.565 82.505 ;
        RECT 115.475 82.035 115.645 82.205 ;
        RECT 115.980 82.035 116.150 82.205 ;
        RECT 116.340 82.035 116.510 82.205 ;
        RECT 114.925 81.855 115.095 82.025 ;
        RECT 117.395 81.975 117.565 82.145 ;
        RECT 114.925 81.495 115.095 81.665 ;
        RECT 115.980 81.605 116.150 81.775 ;
        RECT 116.340 81.605 116.510 81.775 ;
        RECT 117.395 81.615 117.565 81.785 ;
        RECT 114.925 81.135 115.095 81.305 ;
        RECT 115.980 81.175 116.150 81.345 ;
        RECT 116.340 81.175 116.510 81.345 ;
        RECT 116.845 81.175 117.015 81.345 ;
        RECT 117.395 81.255 117.565 81.425 ;
        RECT 114.925 80.775 115.095 80.945 ;
        RECT 115.980 80.745 116.150 80.915 ;
        RECT 116.340 80.745 116.510 80.915 ;
        RECT 117.395 80.895 117.565 81.065 ;
        RECT 117.395 80.535 117.565 80.705 ;
        RECT 114.985 80.115 115.155 80.285 ;
        RECT 115.345 80.115 115.515 80.285 ;
        RECT 115.705 80.115 115.875 80.285 ;
        RECT 116.065 80.115 116.235 80.285 ;
        RECT 116.425 80.115 116.595 80.285 ;
        RECT 116.785 80.115 116.955 80.285 ;
        RECT 117.395 80.175 117.565 80.345 ;
        RECT 118.195 83.660 118.365 83.830 ;
        RECT 118.745 83.720 118.915 83.890 ;
        RECT 119.105 83.720 119.275 83.890 ;
        RECT 119.465 83.720 119.635 83.890 ;
        RECT 119.825 83.720 119.995 83.890 ;
        RECT 120.185 83.720 120.355 83.890 ;
        RECT 120.545 83.720 120.715 83.890 ;
        RECT 120.905 83.720 121.075 83.890 ;
        RECT 118.195 83.300 118.365 83.470 ;
        RECT 118.195 82.940 118.365 83.110 ;
        RECT 119.400 83.090 119.570 83.260 ;
        RECT 119.760 83.090 119.930 83.260 ;
        RECT 120.965 83.200 121.135 83.370 ;
        RECT 120.965 82.840 121.135 83.010 ;
        RECT 118.195 82.580 118.365 82.750 ;
        RECT 118.745 82.660 118.915 82.830 ;
        RECT 119.400 82.660 119.570 82.830 ;
        RECT 119.760 82.660 119.930 82.830 ;
        RECT 120.965 82.480 121.135 82.650 ;
        RECT 118.195 82.220 118.365 82.390 ;
        RECT 119.400 82.230 119.570 82.400 ;
        RECT 119.760 82.230 119.930 82.400 ;
        RECT 118.195 81.860 118.365 82.030 ;
        RECT 120.965 82.120 121.135 82.290 ;
        RECT 118.745 81.800 118.915 81.970 ;
        RECT 119.400 81.800 119.570 81.970 ;
        RECT 119.760 81.800 119.930 81.970 ;
        RECT 118.195 81.500 118.365 81.670 ;
        RECT 120.965 81.760 121.135 81.930 ;
        RECT 119.400 81.370 119.570 81.540 ;
        RECT 119.760 81.370 119.930 81.540 ;
        RECT 120.965 81.400 121.135 81.570 ;
        RECT 118.195 81.140 118.365 81.310 ;
        RECT 118.195 80.780 118.365 80.950 ;
        RECT 118.745 80.940 118.915 81.110 ;
        RECT 119.400 80.940 119.570 81.110 ;
        RECT 119.760 80.940 119.930 81.110 ;
        RECT 120.965 81.040 121.135 81.210 ;
        RECT 120.965 80.680 121.135 80.850 ;
        RECT 118.195 80.420 118.365 80.590 ;
        RECT 119.400 80.510 119.570 80.680 ;
        RECT 119.760 80.510 119.930 80.680 ;
        RECT 120.965 80.320 121.135 80.490 ;
        RECT 109.690 79.720 109.860 79.890 ;
        RECT 110.050 79.720 110.220 79.890 ;
        RECT 111.060 79.720 111.230 79.890 ;
        RECT 111.420 79.720 111.590 79.890 ;
        RECT 112.430 79.720 112.600 79.890 ;
        RECT 112.790 79.720 112.960 79.890 ;
        RECT 108.635 79.540 108.805 79.710 ;
        RECT 113.845 79.710 114.015 79.880 ;
        RECT 108.635 79.180 108.805 79.350 ;
        RECT 108.635 78.820 108.805 78.990 ;
        RECT 108.635 78.460 108.805 78.630 ;
        RECT 71.775 77.890 71.945 78.060 ;
        RECT 72.135 77.890 72.305 78.060 ;
        RECT 72.495 77.890 72.665 78.060 ;
        RECT 72.855 77.890 73.025 78.060 ;
        RECT 73.215 77.890 73.385 78.060 ;
        RECT 73.575 77.890 73.745 78.060 ;
        RECT 75.295 77.890 75.465 78.060 ;
        RECT 75.655 77.890 75.825 78.060 ;
        RECT 76.015 77.890 76.185 78.060 ;
        RECT 76.375 77.890 76.545 78.060 ;
        RECT 76.735 77.890 76.905 78.060 ;
        RECT 77.095 77.890 77.265 78.060 ;
        RECT 77.455 77.890 77.625 78.060 ;
        RECT 77.815 77.890 77.985 78.060 ;
        RECT 78.175 77.890 78.345 78.060 ;
        RECT 78.535 77.890 78.705 78.060 ;
        RECT 78.895 77.890 79.065 78.060 ;
        RECT 79.495 77.890 79.665 78.060 ;
        RECT 79.855 77.890 80.025 78.060 ;
        RECT 80.215 77.890 80.385 78.060 ;
        RECT 80.575 77.890 80.745 78.060 ;
        RECT 80.935 77.890 81.105 78.060 ;
        RECT 81.295 77.890 81.465 78.060 ;
        RECT 81.655 77.890 81.825 78.060 ;
        RECT 82.015 77.890 82.185 78.060 ;
        RECT 82.375 77.890 82.545 78.060 ;
        RECT 82.735 77.890 82.905 78.060 ;
        RECT 83.095 77.890 83.265 78.060 ;
        RECT 84.815 77.890 84.985 78.060 ;
        RECT 85.175 77.890 85.345 78.060 ;
        RECT 85.535 77.890 85.705 78.060 ;
        RECT 85.895 77.890 86.065 78.060 ;
        RECT 86.255 77.890 86.425 78.060 ;
        RECT 86.615 77.890 86.785 78.060 ;
        RECT 108.635 78.100 108.805 78.270 ;
        RECT 108.635 77.740 108.805 77.910 ;
        RECT 110.555 79.300 110.725 79.470 ;
        RECT 110.555 78.940 110.725 79.110 ;
        RECT 110.555 78.580 110.725 78.750 ;
        RECT 110.555 78.220 110.725 78.390 ;
        RECT 110.555 77.860 110.725 78.030 ;
        RECT 111.925 79.300 112.095 79.470 ;
        RECT 111.925 78.940 112.095 79.110 ;
        RECT 111.925 78.580 112.095 78.750 ;
        RECT 111.925 78.220 112.095 78.390 ;
        RECT 111.925 77.860 112.095 78.030 ;
        RECT 113.845 79.350 114.015 79.520 ;
        RECT 118.195 80.060 118.365 80.230 ;
        RECT 119.400 80.080 119.570 80.250 ;
        RECT 119.760 80.080 119.930 80.250 ;
        RECT 120.415 80.080 120.585 80.250 ;
        RECT 120.965 79.960 121.135 80.130 ;
        RECT 119.400 79.650 119.570 79.820 ;
        RECT 119.760 79.650 119.930 79.820 ;
        RECT 113.845 78.990 114.015 79.160 ;
        RECT 113.845 78.630 114.015 78.800 ;
        RECT 113.845 78.270 114.015 78.440 ;
        RECT 113.845 77.910 114.015 78.080 ;
        RECT 108.635 77.380 108.805 77.550 ;
        RECT 109.690 77.440 109.860 77.610 ;
        RECT 110.050 77.440 110.220 77.610 ;
        RECT 111.060 77.440 111.230 77.610 ;
        RECT 111.420 77.440 111.590 77.610 ;
        RECT 112.430 77.440 112.600 77.610 ;
        RECT 112.790 77.440 112.960 77.610 ;
        RECT 113.845 77.550 114.015 77.720 ;
        RECT 113.845 77.190 114.015 77.360 ;
        RECT 108.635 77.020 108.805 77.190 ;
        RECT 108.635 76.660 108.805 76.830 ;
        RECT 108.635 76.300 108.805 76.470 ;
        RECT 108.635 75.940 108.805 76.110 ;
        RECT 108.635 75.580 108.805 75.750 ;
        RECT 110.555 77.020 110.725 77.190 ;
        RECT 110.555 76.660 110.725 76.830 ;
        RECT 110.555 76.300 110.725 76.470 ;
        RECT 110.555 75.940 110.725 76.110 ;
        RECT 110.555 75.580 110.725 75.750 ;
        RECT 111.925 77.020 112.095 77.190 ;
        RECT 111.925 76.660 112.095 76.830 ;
        RECT 111.925 76.300 112.095 76.470 ;
        RECT 111.925 75.940 112.095 76.110 ;
        RECT 111.925 75.580 112.095 75.750 ;
        RECT 113.845 76.830 114.015 77.000 ;
        RECT 113.845 76.470 114.015 76.640 ;
        RECT 113.845 76.110 114.015 76.280 ;
        RECT 113.845 75.750 114.015 75.920 ;
        RECT 108.635 75.220 108.805 75.390 ;
        RECT 113.845 75.390 114.015 75.560 ;
        RECT 114.925 79.265 115.095 79.435 ;
        RECT 115.535 79.325 115.705 79.495 ;
        RECT 115.895 79.325 116.065 79.495 ;
        RECT 116.255 79.325 116.425 79.495 ;
        RECT 116.615 79.325 116.785 79.495 ;
        RECT 116.975 79.325 117.145 79.495 ;
        RECT 117.335 79.325 117.505 79.495 ;
        RECT 114.925 78.905 115.095 79.075 ;
        RECT 114.925 78.545 115.095 78.715 ;
        RECT 115.980 78.655 116.150 78.825 ;
        RECT 116.340 78.655 116.510 78.825 ;
        RECT 117.395 78.705 117.565 78.875 ;
        RECT 114.925 78.185 115.095 78.355 ;
        RECT 115.475 78.225 115.645 78.395 ;
        RECT 115.980 78.225 116.150 78.395 ;
        RECT 116.340 78.225 116.510 78.395 ;
        RECT 117.395 78.345 117.565 78.515 ;
        RECT 114.925 77.825 115.095 77.995 ;
        RECT 117.395 77.985 117.565 78.155 ;
        RECT 115.980 77.795 116.150 77.965 ;
        RECT 116.340 77.795 116.510 77.965 ;
        RECT 117.395 77.625 117.565 77.795 ;
        RECT 115.980 77.365 116.150 77.535 ;
        RECT 116.340 77.365 116.510 77.535 ;
        RECT 116.845 77.365 117.015 77.535 ;
        RECT 114.925 77.185 115.095 77.355 ;
        RECT 117.395 77.265 117.565 77.435 ;
        RECT 114.925 76.825 115.095 76.995 ;
        RECT 115.980 76.935 116.150 77.105 ;
        RECT 116.340 76.935 116.510 77.105 ;
        RECT 117.395 76.905 117.565 77.075 ;
        RECT 114.925 76.465 115.095 76.635 ;
        RECT 115.475 76.505 115.645 76.675 ;
        RECT 115.980 76.505 116.150 76.675 ;
        RECT 116.340 76.505 116.510 76.675 ;
        RECT 117.395 76.545 117.565 76.715 ;
        RECT 114.925 76.105 115.095 76.275 ;
        RECT 115.980 76.075 116.150 76.245 ;
        RECT 116.340 76.075 116.510 76.245 ;
        RECT 117.395 76.185 117.565 76.355 ;
        RECT 117.395 75.825 117.565 75.995 ;
        RECT 114.985 75.405 115.155 75.575 ;
        RECT 115.345 75.405 115.515 75.575 ;
        RECT 115.705 75.405 115.875 75.575 ;
        RECT 116.065 75.405 116.235 75.575 ;
        RECT 116.425 75.405 116.595 75.575 ;
        RECT 116.785 75.405 116.955 75.575 ;
        RECT 117.395 75.465 117.565 75.635 ;
        RECT 118.195 79.470 118.365 79.640 ;
        RECT 120.965 79.600 121.135 79.770 ;
        RECT 118.195 79.110 118.365 79.280 ;
        RECT 119.400 79.220 119.570 79.390 ;
        RECT 119.760 79.220 119.930 79.390 ;
        RECT 120.415 79.220 120.585 79.390 ;
        RECT 120.965 79.240 121.135 79.410 ;
        RECT 118.195 78.750 118.365 78.920 ;
        RECT 119.400 78.790 119.570 78.960 ;
        RECT 119.760 78.790 119.930 78.960 ;
        RECT 120.965 78.880 121.135 79.050 ;
        RECT 118.195 78.390 118.365 78.560 ;
        RECT 118.745 78.360 118.915 78.530 ;
        RECT 119.400 78.360 119.570 78.530 ;
        RECT 119.760 78.360 119.930 78.530 ;
        RECT 120.965 78.520 121.135 78.690 ;
        RECT 118.195 78.030 118.365 78.200 ;
        RECT 120.965 78.160 121.135 78.330 ;
        RECT 119.400 77.930 119.570 78.100 ;
        RECT 119.760 77.930 119.930 78.100 ;
        RECT 118.195 77.670 118.365 77.840 ;
        RECT 120.965 77.800 121.135 77.970 ;
        RECT 118.745 77.500 118.915 77.670 ;
        RECT 119.400 77.500 119.570 77.670 ;
        RECT 119.760 77.500 119.930 77.670 ;
        RECT 118.195 77.310 118.365 77.480 ;
        RECT 120.965 77.440 121.135 77.610 ;
        RECT 118.195 76.950 118.365 77.120 ;
        RECT 119.400 77.070 119.570 77.240 ;
        RECT 119.760 77.070 119.930 77.240 ;
        RECT 120.965 77.080 121.135 77.250 ;
        RECT 118.195 76.590 118.365 76.760 ;
        RECT 118.745 76.640 118.915 76.810 ;
        RECT 119.400 76.640 119.570 76.810 ;
        RECT 119.760 76.640 119.930 76.810 ;
        RECT 120.965 76.720 121.135 76.890 ;
        RECT 121.840 83.860 122.010 84.030 ;
        RECT 121.840 83.500 122.010 83.670 ;
        RECT 121.840 83.140 122.010 83.310 ;
        RECT 121.840 82.780 122.010 82.950 ;
        RECT 121.840 82.420 122.010 82.590 ;
        RECT 122.390 83.860 122.560 84.030 ;
        RECT 122.390 83.500 122.560 83.670 ;
        RECT 122.390 83.140 122.560 83.310 ;
        RECT 122.390 82.780 122.560 82.950 ;
        RECT 122.390 82.420 122.560 82.590 ;
        RECT 125.130 83.860 125.300 84.030 ;
        RECT 125.130 83.500 125.300 83.670 ;
        RECT 125.130 83.140 125.300 83.310 ;
        RECT 125.130 82.780 125.300 82.950 ;
        RECT 125.130 82.420 125.300 82.590 ;
        RECT 125.680 83.710 125.850 83.880 ;
        RECT 125.680 83.350 125.850 83.520 ;
        RECT 125.680 82.990 125.850 83.160 ;
        RECT 125.680 82.630 125.850 82.800 ;
        RECT 121.840 82.060 122.010 82.230 ;
        RECT 125.680 82.270 125.850 82.440 ;
        RECT 122.895 82.000 123.065 82.170 ;
        RECT 123.255 82.000 123.425 82.170 ;
        RECT 124.265 82.000 124.435 82.170 ;
        RECT 124.625 82.000 124.795 82.170 ;
        RECT 121.840 81.700 122.010 81.870 ;
        RECT 125.680 81.910 125.850 82.080 ;
        RECT 121.840 81.340 122.010 81.510 ;
        RECT 121.840 80.980 122.010 81.150 ;
        RECT 121.840 80.620 122.010 80.790 ;
        RECT 121.840 80.260 122.010 80.430 ;
        RECT 122.390 81.580 122.560 81.750 ;
        RECT 122.390 81.220 122.560 81.390 ;
        RECT 122.390 80.860 122.560 81.030 ;
        RECT 122.390 80.500 122.560 80.670 ;
        RECT 122.390 80.140 122.560 80.310 ;
        RECT 125.130 81.580 125.300 81.750 ;
        RECT 125.130 81.220 125.300 81.390 ;
        RECT 125.130 80.860 125.300 81.030 ;
        RECT 125.130 80.500 125.300 80.670 ;
        RECT 125.130 80.140 125.300 80.310 ;
        RECT 125.680 81.550 125.850 81.720 ;
        RECT 125.680 81.190 125.850 81.360 ;
        RECT 125.680 80.830 125.850 81.000 ;
        RECT 125.680 80.470 125.850 80.640 ;
        RECT 121.840 79.900 122.010 80.070 ;
        RECT 125.680 80.110 125.850 80.280 ;
        RECT 122.895 79.720 123.065 79.890 ;
        RECT 123.255 79.720 123.425 79.890 ;
        RECT 124.265 79.720 124.435 79.890 ;
        RECT 124.625 79.720 124.795 79.890 ;
        RECT 125.680 79.750 125.850 79.920 ;
        RECT 121.840 79.540 122.010 79.710 ;
        RECT 121.840 79.180 122.010 79.350 ;
        RECT 121.840 78.820 122.010 78.990 ;
        RECT 121.840 78.460 122.010 78.630 ;
        RECT 121.840 78.100 122.010 78.270 ;
        RECT 121.840 77.740 122.010 77.910 ;
        RECT 122.390 79.300 122.560 79.470 ;
        RECT 122.390 78.940 122.560 79.110 ;
        RECT 122.390 78.580 122.560 78.750 ;
        RECT 122.390 78.220 122.560 78.390 ;
        RECT 122.390 77.860 122.560 78.030 ;
        RECT 123.760 79.300 123.930 79.470 ;
        RECT 123.760 78.940 123.930 79.110 ;
        RECT 123.760 78.580 123.930 78.750 ;
        RECT 123.760 78.220 123.930 78.390 ;
        RECT 123.760 77.860 123.930 78.030 ;
        RECT 125.130 79.300 125.300 79.470 ;
        RECT 125.130 78.940 125.300 79.110 ;
        RECT 125.130 78.580 125.300 78.750 ;
        RECT 125.130 78.220 125.300 78.390 ;
        RECT 125.130 77.860 125.300 78.030 ;
        RECT 125.680 79.390 125.850 79.560 ;
        RECT 125.680 79.030 125.850 79.200 ;
        RECT 125.680 78.670 125.850 78.840 ;
        RECT 125.680 78.310 125.850 78.480 ;
        RECT 125.680 77.950 125.850 78.120 ;
        RECT 121.840 77.380 122.010 77.550 ;
        RECT 122.895 77.440 123.065 77.610 ;
        RECT 123.255 77.440 123.425 77.610 ;
        RECT 124.265 77.440 124.435 77.610 ;
        RECT 124.625 77.440 124.795 77.610 ;
        RECT 125.680 77.590 125.850 77.760 ;
        RECT 125.680 77.230 125.850 77.400 ;
        RECT 121.900 76.810 122.070 76.980 ;
        RECT 122.260 76.810 122.430 76.980 ;
        RECT 122.620 76.810 122.790 76.980 ;
        RECT 122.980 76.810 123.150 76.980 ;
        RECT 123.340 76.810 123.510 76.980 ;
        RECT 123.700 76.810 123.870 76.980 ;
        RECT 124.060 76.810 124.230 76.980 ;
        RECT 124.420 76.810 124.590 76.980 ;
        RECT 124.780 76.810 124.950 76.980 ;
        RECT 125.140 76.810 125.310 76.980 ;
        RECT 125.680 76.870 125.850 77.040 ;
        RECT 118.195 76.230 118.365 76.400 ;
        RECT 119.400 76.210 119.570 76.380 ;
        RECT 119.760 76.210 119.930 76.380 ;
        RECT 120.965 76.360 121.135 76.530 ;
        RECT 120.965 76.000 121.135 76.170 ;
        RECT 118.255 75.580 118.425 75.750 ;
        RECT 118.615 75.580 118.785 75.750 ;
        RECT 118.975 75.580 119.145 75.750 ;
        RECT 119.335 75.580 119.505 75.750 ;
        RECT 119.695 75.580 119.865 75.750 ;
        RECT 120.055 75.580 120.225 75.750 ;
        RECT 120.415 75.580 120.585 75.750 ;
        RECT 120.965 75.640 121.135 75.810 ;
        RECT 109.690 75.160 109.860 75.330 ;
        RECT 110.050 75.160 110.220 75.330 ;
        RECT 111.060 75.160 111.230 75.330 ;
        RECT 111.420 75.160 111.590 75.330 ;
        RECT 112.430 75.160 112.600 75.330 ;
        RECT 112.790 75.160 112.960 75.330 ;
        RECT 108.635 74.860 108.805 75.030 ;
        RECT 113.845 75.030 114.015 75.200 ;
        RECT 108.635 74.500 108.805 74.670 ;
        RECT 108.635 74.140 108.805 74.310 ;
        RECT 108.635 73.780 108.805 73.950 ;
        RECT 108.635 73.420 108.805 73.590 ;
        RECT 110.555 74.740 110.725 74.910 ;
        RECT 110.555 74.380 110.725 74.550 ;
        RECT 110.555 74.020 110.725 74.190 ;
        RECT 110.555 73.660 110.725 73.830 ;
        RECT 110.555 73.300 110.725 73.470 ;
        RECT 111.925 74.740 112.095 74.910 ;
        RECT 111.925 74.380 112.095 74.550 ;
        RECT 111.925 74.020 112.095 74.190 ;
        RECT 111.925 73.660 112.095 73.830 ;
        RECT 111.925 73.300 112.095 73.470 ;
        RECT 113.845 74.670 114.015 74.840 ;
        RECT 113.845 74.310 114.015 74.480 ;
        RECT 113.845 73.950 114.015 74.120 ;
        RECT 113.845 73.590 114.015 73.760 ;
        RECT 108.635 73.060 108.805 73.230 ;
        RECT 113.845 73.230 114.015 73.400 ;
        RECT 109.690 72.880 109.860 73.050 ;
        RECT 110.050 72.880 110.220 73.050 ;
        RECT 111.060 72.880 111.230 73.050 ;
        RECT 111.420 72.880 111.590 73.050 ;
        RECT 112.430 72.880 112.600 73.050 ;
        RECT 112.790 72.880 112.960 73.050 ;
        RECT 108.635 72.700 108.805 72.870 ;
        RECT 65.025 72.360 65.195 72.530 ;
        RECT 65.385 72.360 65.555 72.530 ;
        RECT 65.745 72.360 65.915 72.530 ;
        RECT 66.105 72.360 66.275 72.530 ;
        RECT 66.465 72.360 66.635 72.530 ;
        RECT 66.825 72.360 66.995 72.530 ;
        RECT 68.320 72.360 68.490 72.530 ;
        RECT 68.680 72.360 68.850 72.530 ;
        RECT 69.040 72.360 69.210 72.530 ;
        RECT 69.400 72.360 69.570 72.530 ;
        RECT 69.760 72.360 69.930 72.530 ;
        RECT 70.120 72.360 70.290 72.530 ;
        RECT 70.480 72.360 70.650 72.530 ;
        RECT 70.840 72.360 71.010 72.530 ;
        RECT 64.725 72.010 64.895 72.180 ;
        RECT 71.140 72.010 71.310 72.180 ;
        RECT 64.725 71.650 64.895 71.820 ;
        RECT 65.565 71.690 65.735 71.860 ;
        RECT 65.925 71.690 66.095 71.860 ;
        RECT 68.875 71.690 69.045 71.860 ;
        RECT 69.235 71.690 69.405 71.860 ;
        RECT 69.595 71.690 69.765 71.860 ;
        RECT 69.955 71.690 70.125 71.860 ;
        RECT 70.315 71.690 70.485 71.860 ;
        RECT 71.140 71.650 71.310 71.820 ;
        RECT 64.725 71.290 64.895 71.460 ;
        RECT 66.580 71.440 66.750 71.610 ;
        RECT 65.565 71.260 65.735 71.430 ;
        RECT 65.925 71.260 66.095 71.430 ;
        RECT 64.725 70.930 64.895 71.100 ;
        RECT 66.580 71.080 66.750 71.250 ;
        RECT 68.260 71.440 68.430 71.610 ;
        RECT 68.875 71.260 69.045 71.430 ;
        RECT 69.235 71.260 69.405 71.430 ;
        RECT 69.595 71.260 69.765 71.430 ;
        RECT 69.955 71.260 70.125 71.430 ;
        RECT 70.315 71.260 70.485 71.430 ;
        RECT 71.140 71.290 71.310 71.460 ;
        RECT 68.260 71.080 68.430 71.250 ;
        RECT 65.565 70.830 65.735 71.000 ;
        RECT 65.925 70.830 66.095 71.000 ;
        RECT 68.875 70.830 69.045 71.000 ;
        RECT 69.235 70.830 69.405 71.000 ;
        RECT 69.595 70.830 69.765 71.000 ;
        RECT 69.955 70.830 70.125 71.000 ;
        RECT 70.315 70.830 70.485 71.000 ;
        RECT 71.140 70.930 71.310 71.100 ;
        RECT 64.725 70.570 64.895 70.740 ;
        RECT 66.580 70.580 66.750 70.750 ;
        RECT 65.565 70.400 65.735 70.570 ;
        RECT 65.925 70.400 66.095 70.570 ;
        RECT 64.725 70.210 64.895 70.380 ;
        RECT 66.580 70.220 66.750 70.390 ;
        RECT 68.260 70.580 68.430 70.750 ;
        RECT 71.140 70.570 71.310 70.740 ;
        RECT 68.875 70.400 69.045 70.570 ;
        RECT 69.235 70.400 69.405 70.570 ;
        RECT 69.595 70.400 69.765 70.570 ;
        RECT 69.955 70.400 70.125 70.570 ;
        RECT 70.315 70.400 70.485 70.570 ;
        RECT 68.260 70.220 68.430 70.390 ;
        RECT 71.140 70.210 71.310 70.380 ;
        RECT 64.725 69.850 64.895 70.020 ;
        RECT 65.565 69.970 65.735 70.140 ;
        RECT 65.925 69.970 66.095 70.140 ;
        RECT 68.875 69.970 69.045 70.140 ;
        RECT 69.235 69.970 69.405 70.140 ;
        RECT 69.595 69.970 69.765 70.140 ;
        RECT 69.955 69.970 70.125 70.140 ;
        RECT 70.315 69.970 70.485 70.140 ;
        RECT 66.580 69.720 66.750 69.890 ;
        RECT 64.725 69.490 64.895 69.660 ;
        RECT 65.565 69.540 65.735 69.710 ;
        RECT 65.925 69.540 66.095 69.710 ;
        RECT 66.580 69.360 66.750 69.530 ;
        RECT 68.260 69.720 68.430 69.890 ;
        RECT 71.140 69.850 71.310 70.020 ;
        RECT 68.875 69.540 69.045 69.710 ;
        RECT 69.235 69.540 69.405 69.710 ;
        RECT 69.595 69.540 69.765 69.710 ;
        RECT 69.955 69.540 70.125 69.710 ;
        RECT 70.315 69.540 70.485 69.710 ;
        RECT 68.260 69.360 68.430 69.530 ;
        RECT 71.140 69.490 71.310 69.660 ;
        RECT 64.725 69.130 64.895 69.300 ;
        RECT 65.565 69.110 65.735 69.280 ;
        RECT 65.925 69.110 66.095 69.280 ;
        RECT 68.875 69.110 69.045 69.280 ;
        RECT 69.235 69.110 69.405 69.280 ;
        RECT 69.595 69.110 69.765 69.280 ;
        RECT 69.955 69.110 70.125 69.280 ;
        RECT 70.315 69.110 70.485 69.280 ;
        RECT 71.140 69.130 71.310 69.300 ;
        RECT 64.725 68.770 64.895 68.940 ;
        RECT 66.580 68.860 66.750 69.030 ;
        RECT 65.565 68.680 65.735 68.850 ;
        RECT 65.925 68.680 66.095 68.850 ;
        RECT 64.725 68.410 64.895 68.580 ;
        RECT 66.580 68.500 66.750 68.670 ;
        RECT 68.260 68.860 68.430 69.030 ;
        RECT 68.875 68.680 69.045 68.850 ;
        RECT 69.235 68.680 69.405 68.850 ;
        RECT 69.595 68.680 69.765 68.850 ;
        RECT 69.955 68.680 70.125 68.850 ;
        RECT 70.315 68.680 70.485 68.850 ;
        RECT 71.140 68.770 71.310 68.940 ;
        RECT 68.260 68.500 68.430 68.670 ;
        RECT 65.565 68.250 65.735 68.420 ;
        RECT 65.925 68.250 66.095 68.420 ;
        RECT 68.875 68.250 69.045 68.420 ;
        RECT 69.235 68.250 69.405 68.420 ;
        RECT 69.595 68.250 69.765 68.420 ;
        RECT 69.955 68.250 70.125 68.420 ;
        RECT 70.315 68.250 70.485 68.420 ;
        RECT 71.140 68.410 71.310 68.580 ;
        RECT 64.725 68.050 64.895 68.220 ;
        RECT 66.580 68.000 66.750 68.170 ;
        RECT 64.725 67.690 64.895 67.860 ;
        RECT 65.565 67.820 65.735 67.990 ;
        RECT 65.925 67.820 66.095 67.990 ;
        RECT 66.580 67.640 66.750 67.810 ;
        RECT 68.260 68.000 68.430 68.170 ;
        RECT 71.140 68.050 71.310 68.220 ;
        RECT 68.875 67.820 69.045 67.990 ;
        RECT 69.235 67.820 69.405 67.990 ;
        RECT 69.595 67.820 69.765 67.990 ;
        RECT 69.955 67.820 70.125 67.990 ;
        RECT 70.315 67.820 70.485 67.990 ;
        RECT 68.260 67.640 68.430 67.810 ;
        RECT 71.140 67.690 71.310 67.860 ;
        RECT 64.725 67.330 64.895 67.500 ;
        RECT 65.565 67.390 65.735 67.560 ;
        RECT 65.925 67.390 66.095 67.560 ;
        RECT 68.875 67.390 69.045 67.560 ;
        RECT 69.235 67.390 69.405 67.560 ;
        RECT 69.595 67.390 69.765 67.560 ;
        RECT 69.955 67.390 70.125 67.560 ;
        RECT 70.315 67.390 70.485 67.560 ;
        RECT 71.140 67.330 71.310 67.500 ;
        RECT 64.725 66.970 64.895 67.140 ;
        RECT 66.580 67.140 66.750 67.310 ;
        RECT 65.565 66.960 65.735 67.130 ;
        RECT 65.925 66.960 66.095 67.130 ;
        RECT 66.580 66.780 66.750 66.950 ;
        RECT 68.260 67.140 68.430 67.310 ;
        RECT 68.875 66.960 69.045 67.130 ;
        RECT 69.235 66.960 69.405 67.130 ;
        RECT 69.595 66.960 69.765 67.130 ;
        RECT 69.955 66.960 70.125 67.130 ;
        RECT 70.315 66.960 70.485 67.130 ;
        RECT 71.140 66.970 71.310 67.140 ;
        RECT 68.260 66.780 68.430 66.950 ;
        RECT 64.725 66.610 64.895 66.780 ;
        RECT 65.565 66.530 65.735 66.700 ;
        RECT 65.925 66.530 66.095 66.700 ;
        RECT 68.875 66.530 69.045 66.700 ;
        RECT 69.235 66.530 69.405 66.700 ;
        RECT 69.595 66.530 69.765 66.700 ;
        RECT 69.955 66.530 70.125 66.700 ;
        RECT 70.315 66.530 70.485 66.700 ;
        RECT 71.140 66.610 71.310 66.780 ;
        RECT 64.725 66.250 64.895 66.420 ;
        RECT 66.580 66.280 66.750 66.450 ;
        RECT 65.565 66.100 65.735 66.270 ;
        RECT 65.925 66.100 66.095 66.270 ;
        RECT 64.725 65.890 64.895 66.060 ;
        RECT 66.580 65.920 66.750 66.090 ;
        RECT 68.260 66.280 68.430 66.450 ;
        RECT 68.875 66.100 69.045 66.270 ;
        RECT 69.235 66.100 69.405 66.270 ;
        RECT 69.595 66.100 69.765 66.270 ;
        RECT 69.955 66.100 70.125 66.270 ;
        RECT 70.315 66.100 70.485 66.270 ;
        RECT 71.140 66.250 71.310 66.420 ;
        RECT 68.260 65.920 68.430 66.090 ;
        RECT 71.140 65.890 71.310 66.060 ;
        RECT 64.725 65.530 64.895 65.700 ;
        RECT 65.565 65.670 65.735 65.840 ;
        RECT 65.925 65.670 66.095 65.840 ;
        RECT 68.875 65.670 69.045 65.840 ;
        RECT 69.235 65.670 69.405 65.840 ;
        RECT 69.595 65.670 69.765 65.840 ;
        RECT 69.955 65.670 70.125 65.840 ;
        RECT 70.315 65.670 70.485 65.840 ;
        RECT 66.580 65.420 66.750 65.590 ;
        RECT 64.725 65.170 64.895 65.340 ;
        RECT 65.565 65.240 65.735 65.410 ;
        RECT 65.925 65.240 66.095 65.410 ;
        RECT 66.580 65.060 66.750 65.230 ;
        RECT 68.260 65.420 68.430 65.590 ;
        RECT 71.140 65.530 71.310 65.700 ;
        RECT 68.875 65.240 69.045 65.410 ;
        RECT 69.235 65.240 69.405 65.410 ;
        RECT 69.595 65.240 69.765 65.410 ;
        RECT 69.955 65.240 70.125 65.410 ;
        RECT 70.315 65.240 70.485 65.410 ;
        RECT 68.260 65.060 68.430 65.230 ;
        RECT 71.140 65.170 71.310 65.340 ;
        RECT 64.725 64.810 64.895 64.980 ;
        RECT 65.565 64.810 65.735 64.980 ;
        RECT 65.925 64.810 66.095 64.980 ;
        RECT 68.875 64.810 69.045 64.980 ;
        RECT 69.235 64.810 69.405 64.980 ;
        RECT 69.595 64.810 69.765 64.980 ;
        RECT 69.955 64.810 70.125 64.980 ;
        RECT 70.315 64.810 70.485 64.980 ;
        RECT 71.140 64.810 71.310 64.980 ;
        RECT 64.725 64.450 64.895 64.620 ;
        RECT 66.580 64.560 66.750 64.730 ;
        RECT 65.565 64.380 65.735 64.550 ;
        RECT 65.925 64.380 66.095 64.550 ;
        RECT 64.725 64.090 64.895 64.260 ;
        RECT 66.580 64.200 66.750 64.370 ;
        RECT 68.260 64.560 68.430 64.730 ;
        RECT 68.875 64.380 69.045 64.550 ;
        RECT 69.235 64.380 69.405 64.550 ;
        RECT 69.595 64.380 69.765 64.550 ;
        RECT 69.955 64.380 70.125 64.550 ;
        RECT 70.315 64.380 70.485 64.550 ;
        RECT 71.140 64.450 71.310 64.620 ;
        RECT 68.260 64.200 68.430 64.370 ;
        RECT 65.565 63.950 65.735 64.120 ;
        RECT 65.925 63.950 66.095 64.120 ;
        RECT 68.875 63.950 69.045 64.120 ;
        RECT 69.235 63.950 69.405 64.120 ;
        RECT 69.595 63.950 69.765 64.120 ;
        RECT 69.955 63.950 70.125 64.120 ;
        RECT 70.315 63.950 70.485 64.120 ;
        RECT 71.140 64.090 71.310 64.260 ;
        RECT 64.725 63.730 64.895 63.900 ;
        RECT 71.140 63.730 71.310 63.900 ;
        RECT 65.025 63.280 65.195 63.450 ;
        RECT 65.385 63.280 65.555 63.450 ;
        RECT 65.745 63.280 65.915 63.450 ;
        RECT 66.105 63.280 66.275 63.450 ;
        RECT 66.465 63.280 66.635 63.450 ;
        RECT 66.825 63.280 66.995 63.450 ;
        RECT 68.320 63.280 68.490 63.450 ;
        RECT 68.680 63.280 68.850 63.450 ;
        RECT 69.040 63.280 69.210 63.450 ;
        RECT 69.400 63.280 69.570 63.450 ;
        RECT 69.760 63.280 69.930 63.450 ;
        RECT 70.120 63.280 70.290 63.450 ;
        RECT 70.480 63.280 70.650 63.450 ;
        RECT 70.840 63.280 71.010 63.450 ;
        RECT 74.045 72.360 74.215 72.530 ;
        RECT 74.405 72.360 74.575 72.530 ;
        RECT 74.765 72.360 74.935 72.530 ;
        RECT 75.125 72.360 75.295 72.530 ;
        RECT 75.485 72.360 75.655 72.530 ;
        RECT 75.845 72.360 76.015 72.530 ;
        RECT 77.340 72.360 77.510 72.530 ;
        RECT 77.700 72.360 77.870 72.530 ;
        RECT 78.060 72.360 78.230 72.530 ;
        RECT 78.420 72.360 78.590 72.530 ;
        RECT 78.780 72.360 78.950 72.530 ;
        RECT 79.140 72.360 79.310 72.530 ;
        RECT 79.500 72.360 79.670 72.530 ;
        RECT 79.860 72.360 80.030 72.530 ;
        RECT 80.460 72.360 80.630 72.530 ;
        RECT 80.820 72.360 80.990 72.530 ;
        RECT 81.180 72.360 81.350 72.530 ;
        RECT 81.540 72.360 81.710 72.530 ;
        RECT 81.900 72.360 82.070 72.530 ;
        RECT 82.260 72.360 82.430 72.530 ;
        RECT 82.620 72.360 82.790 72.530 ;
        RECT 82.980 72.360 83.150 72.530 ;
        RECT 84.475 72.360 84.645 72.530 ;
        RECT 84.835 72.360 85.005 72.530 ;
        RECT 85.195 72.360 85.365 72.530 ;
        RECT 85.555 72.360 85.725 72.530 ;
        RECT 85.915 72.360 86.085 72.530 ;
        RECT 86.275 72.360 86.445 72.530 ;
        RECT 73.745 72.010 73.915 72.180 ;
        RECT 80.160 72.010 80.330 72.180 ;
        RECT 73.745 71.650 73.915 71.820 ;
        RECT 74.585 71.690 74.755 71.860 ;
        RECT 74.945 71.690 75.115 71.860 ;
        RECT 77.895 71.690 78.065 71.860 ;
        RECT 78.255 71.690 78.425 71.860 ;
        RECT 78.615 71.690 78.785 71.860 ;
        RECT 78.975 71.690 79.145 71.860 ;
        RECT 79.335 71.690 79.505 71.860 ;
        RECT 86.575 72.010 86.745 72.180 ;
        RECT 80.160 71.650 80.330 71.820 ;
        RECT 80.985 71.690 81.155 71.860 ;
        RECT 81.345 71.690 81.515 71.860 ;
        RECT 81.705 71.690 81.875 71.860 ;
        RECT 82.065 71.690 82.235 71.860 ;
        RECT 82.425 71.690 82.595 71.860 ;
        RECT 85.375 71.690 85.545 71.860 ;
        RECT 85.735 71.690 85.905 71.860 ;
        RECT 73.745 71.290 73.915 71.460 ;
        RECT 75.600 71.440 75.770 71.610 ;
        RECT 74.585 71.260 74.755 71.430 ;
        RECT 74.945 71.260 75.115 71.430 ;
        RECT 73.745 70.930 73.915 71.100 ;
        RECT 75.600 71.080 75.770 71.250 ;
        RECT 77.280 71.440 77.450 71.610 ;
        RECT 86.575 71.650 86.745 71.820 ;
        RECT 77.895 71.260 78.065 71.430 ;
        RECT 78.255 71.260 78.425 71.430 ;
        RECT 78.615 71.260 78.785 71.430 ;
        RECT 78.975 71.260 79.145 71.430 ;
        RECT 79.335 71.260 79.505 71.430 ;
        RECT 80.160 71.290 80.330 71.460 ;
        RECT 83.040 71.440 83.210 71.610 ;
        RECT 77.280 71.080 77.450 71.250 ;
        RECT 80.985 71.260 81.155 71.430 ;
        RECT 81.345 71.260 81.515 71.430 ;
        RECT 81.705 71.260 81.875 71.430 ;
        RECT 82.065 71.260 82.235 71.430 ;
        RECT 82.425 71.260 82.595 71.430 ;
        RECT 74.585 70.830 74.755 71.000 ;
        RECT 74.945 70.830 75.115 71.000 ;
        RECT 77.895 70.830 78.065 71.000 ;
        RECT 78.255 70.830 78.425 71.000 ;
        RECT 78.615 70.830 78.785 71.000 ;
        RECT 78.975 70.830 79.145 71.000 ;
        RECT 79.335 70.830 79.505 71.000 ;
        RECT 80.160 70.930 80.330 71.100 ;
        RECT 83.040 71.080 83.210 71.250 ;
        RECT 84.720 71.440 84.890 71.610 ;
        RECT 85.375 71.260 85.545 71.430 ;
        RECT 85.735 71.260 85.905 71.430 ;
        RECT 86.575 71.290 86.745 71.460 ;
        RECT 84.720 71.080 84.890 71.250 ;
        RECT 73.745 70.570 73.915 70.740 ;
        RECT 75.600 70.580 75.770 70.750 ;
        RECT 74.585 70.400 74.755 70.570 ;
        RECT 74.945 70.400 75.115 70.570 ;
        RECT 73.745 70.210 73.915 70.380 ;
        RECT 75.600 70.220 75.770 70.390 ;
        RECT 77.280 70.580 77.450 70.750 ;
        RECT 80.985 70.830 81.155 71.000 ;
        RECT 81.345 70.830 81.515 71.000 ;
        RECT 81.705 70.830 81.875 71.000 ;
        RECT 82.065 70.830 82.235 71.000 ;
        RECT 82.425 70.830 82.595 71.000 ;
        RECT 85.375 70.830 85.545 71.000 ;
        RECT 85.735 70.830 85.905 71.000 ;
        RECT 86.575 70.930 86.745 71.100 ;
        RECT 80.160 70.570 80.330 70.740 ;
        RECT 83.040 70.580 83.210 70.750 ;
        RECT 77.895 70.400 78.065 70.570 ;
        RECT 78.255 70.400 78.425 70.570 ;
        RECT 78.615 70.400 78.785 70.570 ;
        RECT 78.975 70.400 79.145 70.570 ;
        RECT 79.335 70.400 79.505 70.570 ;
        RECT 77.280 70.220 77.450 70.390 ;
        RECT 80.985 70.400 81.155 70.570 ;
        RECT 81.345 70.400 81.515 70.570 ;
        RECT 81.705 70.400 81.875 70.570 ;
        RECT 82.065 70.400 82.235 70.570 ;
        RECT 82.425 70.400 82.595 70.570 ;
        RECT 80.160 70.210 80.330 70.380 ;
        RECT 83.040 70.220 83.210 70.390 ;
        RECT 84.720 70.580 84.890 70.750 ;
        RECT 86.575 70.570 86.745 70.740 ;
        RECT 85.375 70.400 85.545 70.570 ;
        RECT 85.735 70.400 85.905 70.570 ;
        RECT 84.720 70.220 84.890 70.390 ;
        RECT 73.745 69.850 73.915 70.020 ;
        RECT 74.585 69.970 74.755 70.140 ;
        RECT 74.945 69.970 75.115 70.140 ;
        RECT 77.895 69.970 78.065 70.140 ;
        RECT 78.255 69.970 78.425 70.140 ;
        RECT 78.615 69.970 78.785 70.140 ;
        RECT 78.975 69.970 79.145 70.140 ;
        RECT 79.335 69.970 79.505 70.140 ;
        RECT 86.575 70.210 86.745 70.380 ;
        RECT 75.600 69.720 75.770 69.890 ;
        RECT 73.745 69.490 73.915 69.660 ;
        RECT 74.585 69.540 74.755 69.710 ;
        RECT 74.945 69.540 75.115 69.710 ;
        RECT 75.600 69.360 75.770 69.530 ;
        RECT 77.280 69.720 77.450 69.890 ;
        RECT 80.160 69.850 80.330 70.020 ;
        RECT 80.985 69.970 81.155 70.140 ;
        RECT 81.345 69.970 81.515 70.140 ;
        RECT 81.705 69.970 81.875 70.140 ;
        RECT 82.065 69.970 82.235 70.140 ;
        RECT 82.425 69.970 82.595 70.140 ;
        RECT 85.375 69.970 85.545 70.140 ;
        RECT 85.735 69.970 85.905 70.140 ;
        RECT 77.895 69.540 78.065 69.710 ;
        RECT 78.255 69.540 78.425 69.710 ;
        RECT 78.615 69.540 78.785 69.710 ;
        RECT 78.975 69.540 79.145 69.710 ;
        RECT 79.335 69.540 79.505 69.710 ;
        RECT 83.040 69.720 83.210 69.890 ;
        RECT 77.280 69.360 77.450 69.530 ;
        RECT 80.160 69.490 80.330 69.660 ;
        RECT 80.985 69.540 81.155 69.710 ;
        RECT 81.345 69.540 81.515 69.710 ;
        RECT 81.705 69.540 81.875 69.710 ;
        RECT 82.065 69.540 82.235 69.710 ;
        RECT 82.425 69.540 82.595 69.710 ;
        RECT 73.745 69.130 73.915 69.300 ;
        RECT 83.040 69.360 83.210 69.530 ;
        RECT 84.720 69.720 84.890 69.890 ;
        RECT 86.575 69.850 86.745 70.020 ;
        RECT 85.375 69.540 85.545 69.710 ;
        RECT 85.735 69.540 85.905 69.710 ;
        RECT 84.720 69.360 84.890 69.530 ;
        RECT 86.575 69.490 86.745 69.660 ;
        RECT 74.585 69.110 74.755 69.280 ;
        RECT 74.945 69.110 75.115 69.280 ;
        RECT 77.895 69.110 78.065 69.280 ;
        RECT 78.255 69.110 78.425 69.280 ;
        RECT 78.615 69.110 78.785 69.280 ;
        RECT 78.975 69.110 79.145 69.280 ;
        RECT 79.335 69.110 79.505 69.280 ;
        RECT 80.160 69.130 80.330 69.300 ;
        RECT 73.745 68.770 73.915 68.940 ;
        RECT 75.600 68.860 75.770 69.030 ;
        RECT 74.585 68.680 74.755 68.850 ;
        RECT 74.945 68.680 75.115 68.850 ;
        RECT 73.745 68.410 73.915 68.580 ;
        RECT 75.600 68.500 75.770 68.670 ;
        RECT 77.280 68.860 77.450 69.030 ;
        RECT 80.985 69.110 81.155 69.280 ;
        RECT 81.345 69.110 81.515 69.280 ;
        RECT 81.705 69.110 81.875 69.280 ;
        RECT 82.065 69.110 82.235 69.280 ;
        RECT 82.425 69.110 82.595 69.280 ;
        RECT 85.375 69.110 85.545 69.280 ;
        RECT 85.735 69.110 85.905 69.280 ;
        RECT 86.575 69.130 86.745 69.300 ;
        RECT 77.895 68.680 78.065 68.850 ;
        RECT 78.255 68.680 78.425 68.850 ;
        RECT 78.615 68.680 78.785 68.850 ;
        RECT 78.975 68.680 79.145 68.850 ;
        RECT 79.335 68.680 79.505 68.850 ;
        RECT 80.160 68.770 80.330 68.940 ;
        RECT 83.040 68.860 83.210 69.030 ;
        RECT 77.280 68.500 77.450 68.670 ;
        RECT 80.985 68.680 81.155 68.850 ;
        RECT 81.345 68.680 81.515 68.850 ;
        RECT 81.705 68.680 81.875 68.850 ;
        RECT 82.065 68.680 82.235 68.850 ;
        RECT 82.425 68.680 82.595 68.850 ;
        RECT 74.585 68.250 74.755 68.420 ;
        RECT 74.945 68.250 75.115 68.420 ;
        RECT 77.895 68.250 78.065 68.420 ;
        RECT 78.255 68.250 78.425 68.420 ;
        RECT 78.615 68.250 78.785 68.420 ;
        RECT 78.975 68.250 79.145 68.420 ;
        RECT 79.335 68.250 79.505 68.420 ;
        RECT 80.160 68.410 80.330 68.580 ;
        RECT 83.040 68.500 83.210 68.670 ;
        RECT 84.720 68.860 84.890 69.030 ;
        RECT 85.375 68.680 85.545 68.850 ;
        RECT 85.735 68.680 85.905 68.850 ;
        RECT 86.575 68.770 86.745 68.940 ;
        RECT 84.720 68.500 84.890 68.670 ;
        RECT 73.745 68.050 73.915 68.220 ;
        RECT 80.985 68.250 81.155 68.420 ;
        RECT 81.345 68.250 81.515 68.420 ;
        RECT 81.705 68.250 81.875 68.420 ;
        RECT 82.065 68.250 82.235 68.420 ;
        RECT 82.425 68.250 82.595 68.420 ;
        RECT 85.375 68.250 85.545 68.420 ;
        RECT 85.735 68.250 85.905 68.420 ;
        RECT 86.575 68.410 86.745 68.580 ;
        RECT 75.600 68.000 75.770 68.170 ;
        RECT 73.745 67.690 73.915 67.860 ;
        RECT 74.585 67.820 74.755 67.990 ;
        RECT 74.945 67.820 75.115 67.990 ;
        RECT 75.600 67.640 75.770 67.810 ;
        RECT 77.280 68.000 77.450 68.170 ;
        RECT 80.160 68.050 80.330 68.220 ;
        RECT 77.895 67.820 78.065 67.990 ;
        RECT 78.255 67.820 78.425 67.990 ;
        RECT 78.615 67.820 78.785 67.990 ;
        RECT 78.975 67.820 79.145 67.990 ;
        RECT 79.335 67.820 79.505 67.990 ;
        RECT 83.040 68.000 83.210 68.170 ;
        RECT 77.280 67.640 77.450 67.810 ;
        RECT 80.160 67.690 80.330 67.860 ;
        RECT 80.985 67.820 81.155 67.990 ;
        RECT 81.345 67.820 81.515 67.990 ;
        RECT 81.705 67.820 81.875 67.990 ;
        RECT 82.065 67.820 82.235 67.990 ;
        RECT 82.425 67.820 82.595 67.990 ;
        RECT 73.745 67.330 73.915 67.500 ;
        RECT 74.585 67.390 74.755 67.560 ;
        RECT 74.945 67.390 75.115 67.560 ;
        RECT 77.895 67.390 78.065 67.560 ;
        RECT 78.255 67.390 78.425 67.560 ;
        RECT 78.615 67.390 78.785 67.560 ;
        RECT 78.975 67.390 79.145 67.560 ;
        RECT 79.335 67.390 79.505 67.560 ;
        RECT 83.040 67.640 83.210 67.810 ;
        RECT 84.720 68.000 84.890 68.170 ;
        RECT 86.575 68.050 86.745 68.220 ;
        RECT 85.375 67.820 85.545 67.990 ;
        RECT 85.735 67.820 85.905 67.990 ;
        RECT 84.720 67.640 84.890 67.810 ;
        RECT 86.575 67.690 86.745 67.860 ;
        RECT 80.160 67.330 80.330 67.500 ;
        RECT 80.985 67.390 81.155 67.560 ;
        RECT 81.345 67.390 81.515 67.560 ;
        RECT 81.705 67.390 81.875 67.560 ;
        RECT 82.065 67.390 82.235 67.560 ;
        RECT 82.425 67.390 82.595 67.560 ;
        RECT 85.375 67.390 85.545 67.560 ;
        RECT 85.735 67.390 85.905 67.560 ;
        RECT 73.745 66.970 73.915 67.140 ;
        RECT 75.600 67.140 75.770 67.310 ;
        RECT 74.585 66.960 74.755 67.130 ;
        RECT 74.945 66.960 75.115 67.130 ;
        RECT 75.600 66.780 75.770 66.950 ;
        RECT 77.280 67.140 77.450 67.310 ;
        RECT 86.575 67.330 86.745 67.500 ;
        RECT 77.895 66.960 78.065 67.130 ;
        RECT 78.255 66.960 78.425 67.130 ;
        RECT 78.615 66.960 78.785 67.130 ;
        RECT 78.975 66.960 79.145 67.130 ;
        RECT 79.335 66.960 79.505 67.130 ;
        RECT 80.160 66.970 80.330 67.140 ;
        RECT 83.040 67.140 83.210 67.310 ;
        RECT 77.280 66.780 77.450 66.950 ;
        RECT 80.985 66.960 81.155 67.130 ;
        RECT 81.345 66.960 81.515 67.130 ;
        RECT 81.705 66.960 81.875 67.130 ;
        RECT 82.065 66.960 82.235 67.130 ;
        RECT 82.425 66.960 82.595 67.130 ;
        RECT 83.040 66.780 83.210 66.950 ;
        RECT 84.720 67.140 84.890 67.310 ;
        RECT 85.375 66.960 85.545 67.130 ;
        RECT 85.735 66.960 85.905 67.130 ;
        RECT 86.575 66.970 86.745 67.140 ;
        RECT 84.720 66.780 84.890 66.950 ;
        RECT 73.745 66.610 73.915 66.780 ;
        RECT 74.585 66.530 74.755 66.700 ;
        RECT 74.945 66.530 75.115 66.700 ;
        RECT 77.895 66.530 78.065 66.700 ;
        RECT 78.255 66.530 78.425 66.700 ;
        RECT 78.615 66.530 78.785 66.700 ;
        RECT 78.975 66.530 79.145 66.700 ;
        RECT 79.335 66.530 79.505 66.700 ;
        RECT 80.160 66.610 80.330 66.780 ;
        RECT 73.745 66.250 73.915 66.420 ;
        RECT 75.600 66.280 75.770 66.450 ;
        RECT 74.585 66.100 74.755 66.270 ;
        RECT 74.945 66.100 75.115 66.270 ;
        RECT 73.745 65.890 73.915 66.060 ;
        RECT 75.600 65.920 75.770 66.090 ;
        RECT 77.280 66.280 77.450 66.450 ;
        RECT 80.985 66.530 81.155 66.700 ;
        RECT 81.345 66.530 81.515 66.700 ;
        RECT 81.705 66.530 81.875 66.700 ;
        RECT 82.065 66.530 82.235 66.700 ;
        RECT 82.425 66.530 82.595 66.700 ;
        RECT 85.375 66.530 85.545 66.700 ;
        RECT 85.735 66.530 85.905 66.700 ;
        RECT 86.575 66.610 86.745 66.780 ;
        RECT 77.895 66.100 78.065 66.270 ;
        RECT 78.255 66.100 78.425 66.270 ;
        RECT 78.615 66.100 78.785 66.270 ;
        RECT 78.975 66.100 79.145 66.270 ;
        RECT 79.335 66.100 79.505 66.270 ;
        RECT 80.160 66.250 80.330 66.420 ;
        RECT 83.040 66.280 83.210 66.450 ;
        RECT 77.280 65.920 77.450 66.090 ;
        RECT 80.985 66.100 81.155 66.270 ;
        RECT 81.345 66.100 81.515 66.270 ;
        RECT 81.705 66.100 81.875 66.270 ;
        RECT 82.065 66.100 82.235 66.270 ;
        RECT 82.425 66.100 82.595 66.270 ;
        RECT 80.160 65.890 80.330 66.060 ;
        RECT 83.040 65.920 83.210 66.090 ;
        RECT 84.720 66.280 84.890 66.450 ;
        RECT 85.375 66.100 85.545 66.270 ;
        RECT 85.735 66.100 85.905 66.270 ;
        RECT 86.575 66.250 86.745 66.420 ;
        RECT 84.720 65.920 84.890 66.090 ;
        RECT 73.745 65.530 73.915 65.700 ;
        RECT 74.585 65.670 74.755 65.840 ;
        RECT 74.945 65.670 75.115 65.840 ;
        RECT 77.895 65.670 78.065 65.840 ;
        RECT 78.255 65.670 78.425 65.840 ;
        RECT 78.615 65.670 78.785 65.840 ;
        RECT 78.975 65.670 79.145 65.840 ;
        RECT 79.335 65.670 79.505 65.840 ;
        RECT 86.575 65.890 86.745 66.060 ;
        RECT 75.600 65.420 75.770 65.590 ;
        RECT 73.745 65.170 73.915 65.340 ;
        RECT 74.585 65.240 74.755 65.410 ;
        RECT 74.945 65.240 75.115 65.410 ;
        RECT 75.600 65.060 75.770 65.230 ;
        RECT 77.280 65.420 77.450 65.590 ;
        RECT 80.160 65.530 80.330 65.700 ;
        RECT 80.985 65.670 81.155 65.840 ;
        RECT 81.345 65.670 81.515 65.840 ;
        RECT 81.705 65.670 81.875 65.840 ;
        RECT 82.065 65.670 82.235 65.840 ;
        RECT 82.425 65.670 82.595 65.840 ;
        RECT 85.375 65.670 85.545 65.840 ;
        RECT 85.735 65.670 85.905 65.840 ;
        RECT 77.895 65.240 78.065 65.410 ;
        RECT 78.255 65.240 78.425 65.410 ;
        RECT 78.615 65.240 78.785 65.410 ;
        RECT 78.975 65.240 79.145 65.410 ;
        RECT 79.335 65.240 79.505 65.410 ;
        RECT 83.040 65.420 83.210 65.590 ;
        RECT 77.280 65.060 77.450 65.230 ;
        RECT 80.160 65.170 80.330 65.340 ;
        RECT 80.985 65.240 81.155 65.410 ;
        RECT 81.345 65.240 81.515 65.410 ;
        RECT 81.705 65.240 81.875 65.410 ;
        RECT 82.065 65.240 82.235 65.410 ;
        RECT 82.425 65.240 82.595 65.410 ;
        RECT 83.040 65.060 83.210 65.230 ;
        RECT 84.720 65.420 84.890 65.590 ;
        RECT 86.575 65.530 86.745 65.700 ;
        RECT 85.375 65.240 85.545 65.410 ;
        RECT 85.735 65.240 85.905 65.410 ;
        RECT 84.720 65.060 84.890 65.230 ;
        RECT 86.575 65.170 86.745 65.340 ;
        RECT 73.745 64.810 73.915 64.980 ;
        RECT 74.585 64.810 74.755 64.980 ;
        RECT 74.945 64.810 75.115 64.980 ;
        RECT 77.895 64.810 78.065 64.980 ;
        RECT 78.255 64.810 78.425 64.980 ;
        RECT 78.615 64.810 78.785 64.980 ;
        RECT 78.975 64.810 79.145 64.980 ;
        RECT 79.335 64.810 79.505 64.980 ;
        RECT 80.160 64.810 80.330 64.980 ;
        RECT 80.985 64.810 81.155 64.980 ;
        RECT 81.345 64.810 81.515 64.980 ;
        RECT 81.705 64.810 81.875 64.980 ;
        RECT 82.065 64.810 82.235 64.980 ;
        RECT 82.425 64.810 82.595 64.980 ;
        RECT 85.375 64.810 85.545 64.980 ;
        RECT 85.735 64.810 85.905 64.980 ;
        RECT 86.575 64.810 86.745 64.980 ;
        RECT 73.745 64.450 73.915 64.620 ;
        RECT 75.600 64.560 75.770 64.730 ;
        RECT 74.585 64.380 74.755 64.550 ;
        RECT 74.945 64.380 75.115 64.550 ;
        RECT 73.745 64.090 73.915 64.260 ;
        RECT 75.600 64.200 75.770 64.370 ;
        RECT 77.280 64.560 77.450 64.730 ;
        RECT 77.895 64.380 78.065 64.550 ;
        RECT 78.255 64.380 78.425 64.550 ;
        RECT 78.615 64.380 78.785 64.550 ;
        RECT 78.975 64.380 79.145 64.550 ;
        RECT 79.335 64.380 79.505 64.550 ;
        RECT 80.160 64.450 80.330 64.620 ;
        RECT 83.040 64.560 83.210 64.730 ;
        RECT 77.280 64.200 77.450 64.370 ;
        RECT 80.985 64.380 81.155 64.550 ;
        RECT 81.345 64.380 81.515 64.550 ;
        RECT 81.705 64.380 81.875 64.550 ;
        RECT 82.065 64.380 82.235 64.550 ;
        RECT 82.425 64.380 82.595 64.550 ;
        RECT 74.585 63.950 74.755 64.120 ;
        RECT 74.945 63.950 75.115 64.120 ;
        RECT 77.895 63.950 78.065 64.120 ;
        RECT 78.255 63.950 78.425 64.120 ;
        RECT 78.615 63.950 78.785 64.120 ;
        RECT 78.975 63.950 79.145 64.120 ;
        RECT 79.335 63.950 79.505 64.120 ;
        RECT 80.160 64.090 80.330 64.260 ;
        RECT 83.040 64.200 83.210 64.370 ;
        RECT 84.720 64.560 84.890 64.730 ;
        RECT 85.375 64.380 85.545 64.550 ;
        RECT 85.735 64.380 85.905 64.550 ;
        RECT 86.575 64.450 86.745 64.620 ;
        RECT 84.720 64.200 84.890 64.370 ;
        RECT 73.745 63.730 73.915 63.900 ;
        RECT 80.985 63.950 81.155 64.120 ;
        RECT 81.345 63.950 81.515 64.120 ;
        RECT 81.705 63.950 81.875 64.120 ;
        RECT 82.065 63.950 82.235 64.120 ;
        RECT 82.425 63.950 82.595 64.120 ;
        RECT 85.375 63.950 85.545 64.120 ;
        RECT 85.735 63.950 85.905 64.120 ;
        RECT 86.575 64.090 86.745 64.260 ;
        RECT 80.160 63.730 80.330 63.900 ;
        RECT 86.575 63.730 86.745 63.900 ;
        RECT 74.045 63.280 74.215 63.450 ;
        RECT 74.405 63.280 74.575 63.450 ;
        RECT 74.765 63.280 74.935 63.450 ;
        RECT 75.125 63.280 75.295 63.450 ;
        RECT 75.485 63.280 75.655 63.450 ;
        RECT 75.845 63.280 76.015 63.450 ;
        RECT 77.340 63.280 77.510 63.450 ;
        RECT 77.700 63.280 77.870 63.450 ;
        RECT 78.060 63.280 78.230 63.450 ;
        RECT 78.420 63.280 78.590 63.450 ;
        RECT 78.780 63.280 78.950 63.450 ;
        RECT 79.140 63.280 79.310 63.450 ;
        RECT 79.500 63.280 79.670 63.450 ;
        RECT 79.860 63.280 80.030 63.450 ;
        RECT 80.460 63.280 80.630 63.450 ;
        RECT 80.820 63.280 80.990 63.450 ;
        RECT 81.180 63.280 81.350 63.450 ;
        RECT 81.540 63.280 81.710 63.450 ;
        RECT 81.900 63.280 82.070 63.450 ;
        RECT 82.260 63.280 82.430 63.450 ;
        RECT 82.620 63.280 82.790 63.450 ;
        RECT 82.980 63.280 83.150 63.450 ;
        RECT 84.475 63.280 84.645 63.450 ;
        RECT 84.835 63.280 85.005 63.450 ;
        RECT 85.195 63.280 85.365 63.450 ;
        RECT 85.555 63.280 85.725 63.450 ;
        RECT 85.915 63.280 86.085 63.450 ;
        RECT 86.275 63.280 86.445 63.450 ;
        RECT 88.805 72.360 88.975 72.530 ;
        RECT 89.165 72.360 89.335 72.530 ;
        RECT 89.525 72.360 89.695 72.530 ;
        RECT 89.885 72.360 90.055 72.530 ;
        RECT 90.245 72.360 90.415 72.530 ;
        RECT 90.605 72.360 90.775 72.530 ;
        RECT 92.100 72.360 92.270 72.530 ;
        RECT 92.460 72.360 92.630 72.530 ;
        RECT 92.820 72.360 92.990 72.530 ;
        RECT 93.180 72.360 93.350 72.530 ;
        RECT 93.540 72.360 93.710 72.530 ;
        RECT 93.900 72.360 94.070 72.530 ;
        RECT 94.260 72.360 94.430 72.530 ;
        RECT 94.620 72.360 94.790 72.530 ;
        RECT 88.505 72.010 88.675 72.180 ;
        RECT 94.920 72.010 95.090 72.180 ;
        RECT 88.505 71.650 88.675 71.820 ;
        RECT 89.345 71.690 89.515 71.860 ;
        RECT 89.705 71.690 89.875 71.860 ;
        RECT 92.655 71.690 92.825 71.860 ;
        RECT 93.015 71.690 93.185 71.860 ;
        RECT 93.375 71.690 93.545 71.860 ;
        RECT 93.735 71.690 93.905 71.860 ;
        RECT 94.095 71.690 94.265 71.860 ;
        RECT 94.920 71.650 95.090 71.820 ;
        RECT 88.505 71.290 88.675 71.460 ;
        RECT 90.360 71.440 90.530 71.610 ;
        RECT 89.345 71.260 89.515 71.430 ;
        RECT 89.705 71.260 89.875 71.430 ;
        RECT 88.505 70.930 88.675 71.100 ;
        RECT 90.360 71.080 90.530 71.250 ;
        RECT 92.040 71.440 92.210 71.610 ;
        RECT 92.655 71.260 92.825 71.430 ;
        RECT 93.015 71.260 93.185 71.430 ;
        RECT 93.375 71.260 93.545 71.430 ;
        RECT 93.735 71.260 93.905 71.430 ;
        RECT 94.095 71.260 94.265 71.430 ;
        RECT 94.920 71.290 95.090 71.460 ;
        RECT 92.040 71.080 92.210 71.250 ;
        RECT 89.345 70.830 89.515 71.000 ;
        RECT 89.705 70.830 89.875 71.000 ;
        RECT 92.655 70.830 92.825 71.000 ;
        RECT 93.015 70.830 93.185 71.000 ;
        RECT 93.375 70.830 93.545 71.000 ;
        RECT 93.735 70.830 93.905 71.000 ;
        RECT 94.095 70.830 94.265 71.000 ;
        RECT 94.920 70.930 95.090 71.100 ;
        RECT 88.505 70.570 88.675 70.740 ;
        RECT 90.360 70.580 90.530 70.750 ;
        RECT 89.345 70.400 89.515 70.570 ;
        RECT 89.705 70.400 89.875 70.570 ;
        RECT 88.505 70.210 88.675 70.380 ;
        RECT 90.360 70.220 90.530 70.390 ;
        RECT 92.040 70.580 92.210 70.750 ;
        RECT 94.920 70.570 95.090 70.740 ;
        RECT 92.655 70.400 92.825 70.570 ;
        RECT 93.015 70.400 93.185 70.570 ;
        RECT 93.375 70.400 93.545 70.570 ;
        RECT 93.735 70.400 93.905 70.570 ;
        RECT 94.095 70.400 94.265 70.570 ;
        RECT 92.040 70.220 92.210 70.390 ;
        RECT 94.920 70.210 95.090 70.380 ;
        RECT 88.505 69.850 88.675 70.020 ;
        RECT 89.345 69.970 89.515 70.140 ;
        RECT 89.705 69.970 89.875 70.140 ;
        RECT 92.655 69.970 92.825 70.140 ;
        RECT 93.015 69.970 93.185 70.140 ;
        RECT 93.375 69.970 93.545 70.140 ;
        RECT 93.735 69.970 93.905 70.140 ;
        RECT 94.095 69.970 94.265 70.140 ;
        RECT 90.360 69.720 90.530 69.890 ;
        RECT 88.505 69.490 88.675 69.660 ;
        RECT 89.345 69.540 89.515 69.710 ;
        RECT 89.705 69.540 89.875 69.710 ;
        RECT 90.360 69.360 90.530 69.530 ;
        RECT 92.040 69.720 92.210 69.890 ;
        RECT 94.920 69.850 95.090 70.020 ;
        RECT 92.655 69.540 92.825 69.710 ;
        RECT 93.015 69.540 93.185 69.710 ;
        RECT 93.375 69.540 93.545 69.710 ;
        RECT 93.735 69.540 93.905 69.710 ;
        RECT 94.095 69.540 94.265 69.710 ;
        RECT 92.040 69.360 92.210 69.530 ;
        RECT 94.920 69.490 95.090 69.660 ;
        RECT 88.505 69.130 88.675 69.300 ;
        RECT 89.345 69.110 89.515 69.280 ;
        RECT 89.705 69.110 89.875 69.280 ;
        RECT 92.655 69.110 92.825 69.280 ;
        RECT 93.015 69.110 93.185 69.280 ;
        RECT 93.375 69.110 93.545 69.280 ;
        RECT 93.735 69.110 93.905 69.280 ;
        RECT 94.095 69.110 94.265 69.280 ;
        RECT 94.920 69.130 95.090 69.300 ;
        RECT 88.505 68.770 88.675 68.940 ;
        RECT 90.360 68.860 90.530 69.030 ;
        RECT 89.345 68.680 89.515 68.850 ;
        RECT 89.705 68.680 89.875 68.850 ;
        RECT 88.505 68.410 88.675 68.580 ;
        RECT 90.360 68.500 90.530 68.670 ;
        RECT 92.040 68.860 92.210 69.030 ;
        RECT 92.655 68.680 92.825 68.850 ;
        RECT 93.015 68.680 93.185 68.850 ;
        RECT 93.375 68.680 93.545 68.850 ;
        RECT 93.735 68.680 93.905 68.850 ;
        RECT 94.095 68.680 94.265 68.850 ;
        RECT 94.920 68.770 95.090 68.940 ;
        RECT 92.040 68.500 92.210 68.670 ;
        RECT 89.345 68.250 89.515 68.420 ;
        RECT 89.705 68.250 89.875 68.420 ;
        RECT 92.655 68.250 92.825 68.420 ;
        RECT 93.015 68.250 93.185 68.420 ;
        RECT 93.375 68.250 93.545 68.420 ;
        RECT 93.735 68.250 93.905 68.420 ;
        RECT 94.095 68.250 94.265 68.420 ;
        RECT 94.920 68.410 95.090 68.580 ;
        RECT 88.505 68.050 88.675 68.220 ;
        RECT 90.360 68.000 90.530 68.170 ;
        RECT 88.505 67.690 88.675 67.860 ;
        RECT 89.345 67.820 89.515 67.990 ;
        RECT 89.705 67.820 89.875 67.990 ;
        RECT 90.360 67.640 90.530 67.810 ;
        RECT 92.040 68.000 92.210 68.170 ;
        RECT 94.920 68.050 95.090 68.220 ;
        RECT 92.655 67.820 92.825 67.990 ;
        RECT 93.015 67.820 93.185 67.990 ;
        RECT 93.375 67.820 93.545 67.990 ;
        RECT 93.735 67.820 93.905 67.990 ;
        RECT 94.095 67.820 94.265 67.990 ;
        RECT 92.040 67.640 92.210 67.810 ;
        RECT 94.920 67.690 95.090 67.860 ;
        RECT 88.505 67.330 88.675 67.500 ;
        RECT 89.345 67.390 89.515 67.560 ;
        RECT 89.705 67.390 89.875 67.560 ;
        RECT 92.655 67.390 92.825 67.560 ;
        RECT 93.015 67.390 93.185 67.560 ;
        RECT 93.375 67.390 93.545 67.560 ;
        RECT 93.735 67.390 93.905 67.560 ;
        RECT 94.095 67.390 94.265 67.560 ;
        RECT 94.920 67.330 95.090 67.500 ;
        RECT 88.505 66.970 88.675 67.140 ;
        RECT 90.360 67.140 90.530 67.310 ;
        RECT 89.345 66.960 89.515 67.130 ;
        RECT 89.705 66.960 89.875 67.130 ;
        RECT 90.360 66.780 90.530 66.950 ;
        RECT 92.040 67.140 92.210 67.310 ;
        RECT 92.655 66.960 92.825 67.130 ;
        RECT 93.015 66.960 93.185 67.130 ;
        RECT 93.375 66.960 93.545 67.130 ;
        RECT 93.735 66.960 93.905 67.130 ;
        RECT 94.095 66.960 94.265 67.130 ;
        RECT 94.920 66.970 95.090 67.140 ;
        RECT 92.040 66.780 92.210 66.950 ;
        RECT 88.505 66.610 88.675 66.780 ;
        RECT 89.345 66.530 89.515 66.700 ;
        RECT 89.705 66.530 89.875 66.700 ;
        RECT 92.655 66.530 92.825 66.700 ;
        RECT 93.015 66.530 93.185 66.700 ;
        RECT 93.375 66.530 93.545 66.700 ;
        RECT 93.735 66.530 93.905 66.700 ;
        RECT 94.095 66.530 94.265 66.700 ;
        RECT 94.920 66.610 95.090 66.780 ;
        RECT 88.505 66.250 88.675 66.420 ;
        RECT 90.360 66.280 90.530 66.450 ;
        RECT 89.345 66.100 89.515 66.270 ;
        RECT 89.705 66.100 89.875 66.270 ;
        RECT 88.505 65.890 88.675 66.060 ;
        RECT 90.360 65.920 90.530 66.090 ;
        RECT 92.040 66.280 92.210 66.450 ;
        RECT 92.655 66.100 92.825 66.270 ;
        RECT 93.015 66.100 93.185 66.270 ;
        RECT 93.375 66.100 93.545 66.270 ;
        RECT 93.735 66.100 93.905 66.270 ;
        RECT 94.095 66.100 94.265 66.270 ;
        RECT 94.920 66.250 95.090 66.420 ;
        RECT 92.040 65.920 92.210 66.090 ;
        RECT 94.920 65.890 95.090 66.060 ;
        RECT 88.505 65.530 88.675 65.700 ;
        RECT 89.345 65.670 89.515 65.840 ;
        RECT 89.705 65.670 89.875 65.840 ;
        RECT 92.655 65.670 92.825 65.840 ;
        RECT 93.015 65.670 93.185 65.840 ;
        RECT 93.375 65.670 93.545 65.840 ;
        RECT 93.735 65.670 93.905 65.840 ;
        RECT 94.095 65.670 94.265 65.840 ;
        RECT 90.360 65.420 90.530 65.590 ;
        RECT 88.505 65.170 88.675 65.340 ;
        RECT 89.345 65.240 89.515 65.410 ;
        RECT 89.705 65.240 89.875 65.410 ;
        RECT 90.360 65.060 90.530 65.230 ;
        RECT 92.040 65.420 92.210 65.590 ;
        RECT 94.920 65.530 95.090 65.700 ;
        RECT 92.655 65.240 92.825 65.410 ;
        RECT 93.015 65.240 93.185 65.410 ;
        RECT 93.375 65.240 93.545 65.410 ;
        RECT 93.735 65.240 93.905 65.410 ;
        RECT 94.095 65.240 94.265 65.410 ;
        RECT 92.040 65.060 92.210 65.230 ;
        RECT 94.920 65.170 95.090 65.340 ;
        RECT 88.505 64.810 88.675 64.980 ;
        RECT 89.345 64.810 89.515 64.980 ;
        RECT 89.705 64.810 89.875 64.980 ;
        RECT 92.655 64.810 92.825 64.980 ;
        RECT 93.015 64.810 93.185 64.980 ;
        RECT 93.375 64.810 93.545 64.980 ;
        RECT 93.735 64.810 93.905 64.980 ;
        RECT 94.095 64.810 94.265 64.980 ;
        RECT 94.920 64.810 95.090 64.980 ;
        RECT 88.505 64.450 88.675 64.620 ;
        RECT 90.360 64.560 90.530 64.730 ;
        RECT 89.345 64.380 89.515 64.550 ;
        RECT 89.705 64.380 89.875 64.550 ;
        RECT 88.505 64.090 88.675 64.260 ;
        RECT 90.360 64.200 90.530 64.370 ;
        RECT 92.040 64.560 92.210 64.730 ;
        RECT 92.655 64.380 92.825 64.550 ;
        RECT 93.015 64.380 93.185 64.550 ;
        RECT 93.375 64.380 93.545 64.550 ;
        RECT 93.735 64.380 93.905 64.550 ;
        RECT 94.095 64.380 94.265 64.550 ;
        RECT 94.920 64.450 95.090 64.620 ;
        RECT 92.040 64.200 92.210 64.370 ;
        RECT 89.345 63.950 89.515 64.120 ;
        RECT 89.705 63.950 89.875 64.120 ;
        RECT 92.655 63.950 92.825 64.120 ;
        RECT 93.015 63.950 93.185 64.120 ;
        RECT 93.375 63.950 93.545 64.120 ;
        RECT 93.735 63.950 93.905 64.120 ;
        RECT 94.095 63.950 94.265 64.120 ;
        RECT 94.920 64.090 95.090 64.260 ;
        RECT 88.505 63.730 88.675 63.900 ;
        RECT 94.920 63.730 95.090 63.900 ;
        RECT 88.805 63.280 88.975 63.450 ;
        RECT 89.165 63.280 89.335 63.450 ;
        RECT 89.525 63.280 89.695 63.450 ;
        RECT 89.885 63.280 90.055 63.450 ;
        RECT 90.245 63.280 90.415 63.450 ;
        RECT 90.605 63.280 90.775 63.450 ;
        RECT 92.100 63.280 92.270 63.450 ;
        RECT 92.460 63.280 92.630 63.450 ;
        RECT 92.820 63.280 92.990 63.450 ;
        RECT 93.180 63.280 93.350 63.450 ;
        RECT 93.540 63.280 93.710 63.450 ;
        RECT 93.900 63.280 94.070 63.450 ;
        RECT 94.260 63.280 94.430 63.450 ;
        RECT 94.620 63.280 94.790 63.450 ;
        RECT 113.845 72.870 114.015 73.040 ;
        RECT 108.635 72.340 108.805 72.510 ;
        RECT 108.635 71.980 108.805 72.150 ;
        RECT 108.635 71.620 108.805 71.790 ;
        RECT 108.635 71.260 108.805 71.430 ;
        RECT 108.635 70.900 108.805 71.070 ;
        RECT 110.555 72.460 110.725 72.630 ;
        RECT 110.555 72.100 110.725 72.270 ;
        RECT 110.555 71.740 110.725 71.910 ;
        RECT 110.555 71.380 110.725 71.550 ;
        RECT 110.555 71.020 110.725 71.190 ;
        RECT 111.925 72.460 112.095 72.630 ;
        RECT 111.925 72.100 112.095 72.270 ;
        RECT 111.925 71.740 112.095 71.910 ;
        RECT 111.925 71.380 112.095 71.550 ;
        RECT 111.925 71.020 112.095 71.190 ;
        RECT 113.845 72.510 114.015 72.680 ;
        RECT 113.845 72.150 114.015 72.320 ;
        RECT 113.845 71.790 114.015 71.960 ;
        RECT 113.845 71.430 114.015 71.600 ;
        RECT 113.845 71.070 114.015 71.240 ;
        RECT 108.635 70.540 108.805 70.710 ;
        RECT 109.690 70.600 109.860 70.770 ;
        RECT 110.050 70.600 110.220 70.770 ;
        RECT 111.060 70.600 111.230 70.770 ;
        RECT 111.420 70.600 111.590 70.770 ;
        RECT 112.430 70.600 112.600 70.770 ;
        RECT 112.790 70.600 112.960 70.770 ;
        RECT 113.845 70.710 114.015 70.880 ;
        RECT 113.845 70.350 114.015 70.520 ;
        RECT 108.635 70.180 108.805 70.350 ;
        RECT 108.635 69.820 108.805 69.990 ;
        RECT 108.635 69.460 108.805 69.630 ;
        RECT 108.635 69.100 108.805 69.270 ;
        RECT 108.635 68.740 108.805 68.910 ;
        RECT 110.555 70.180 110.725 70.350 ;
        RECT 110.555 69.820 110.725 69.990 ;
        RECT 110.555 69.460 110.725 69.630 ;
        RECT 110.555 69.100 110.725 69.270 ;
        RECT 110.555 68.740 110.725 68.910 ;
        RECT 111.925 70.180 112.095 70.350 ;
        RECT 111.925 69.820 112.095 69.990 ;
        RECT 111.925 69.460 112.095 69.630 ;
        RECT 111.925 69.100 112.095 69.270 ;
        RECT 111.925 68.740 112.095 68.910 ;
        RECT 113.845 69.990 114.015 70.160 ;
        RECT 113.845 69.630 114.015 69.800 ;
        RECT 113.845 69.270 114.015 69.440 ;
        RECT 113.845 68.910 114.015 69.080 ;
        RECT 108.635 68.380 108.805 68.550 ;
        RECT 113.845 68.550 114.015 68.720 ;
        RECT 109.690 68.320 109.860 68.490 ;
        RECT 110.050 68.320 110.220 68.490 ;
        RECT 111.060 68.320 111.230 68.490 ;
        RECT 111.420 68.320 111.590 68.490 ;
        RECT 112.430 68.320 112.600 68.490 ;
        RECT 112.790 68.320 112.960 68.490 ;
        RECT 108.635 68.020 108.805 68.190 ;
        RECT 113.845 68.190 114.015 68.360 ;
        RECT 108.635 67.660 108.805 67.830 ;
        RECT 108.635 67.300 108.805 67.470 ;
        RECT 108.635 66.940 108.805 67.110 ;
        RECT 108.635 66.580 108.805 66.750 ;
        RECT 110.555 67.900 110.725 68.070 ;
        RECT 110.555 67.540 110.725 67.710 ;
        RECT 110.555 67.180 110.725 67.350 ;
        RECT 110.555 66.820 110.725 66.990 ;
        RECT 110.555 66.460 110.725 66.630 ;
        RECT 111.925 67.900 112.095 68.070 ;
        RECT 111.925 67.540 112.095 67.710 ;
        RECT 111.925 67.180 112.095 67.350 ;
        RECT 111.925 66.820 112.095 66.990 ;
        RECT 111.925 66.460 112.095 66.630 ;
        RECT 113.845 67.830 114.015 68.000 ;
        RECT 113.845 67.470 114.015 67.640 ;
        RECT 113.845 67.110 114.015 67.280 ;
        RECT 113.845 66.750 114.015 66.920 ;
        RECT 108.635 66.220 108.805 66.390 ;
        RECT 113.845 66.390 114.015 66.560 ;
        RECT 109.690 66.040 109.860 66.210 ;
        RECT 110.050 66.040 110.220 66.210 ;
        RECT 111.060 66.040 111.230 66.210 ;
        RECT 111.420 66.040 111.590 66.210 ;
        RECT 112.430 66.040 112.600 66.210 ;
        RECT 112.790 66.040 112.960 66.210 ;
        RECT 108.635 65.860 108.805 66.030 ;
        RECT 113.845 66.030 114.015 66.200 ;
        RECT 108.635 65.500 108.805 65.670 ;
        RECT 108.635 65.140 108.805 65.310 ;
        RECT 108.635 64.780 108.805 64.950 ;
        RECT 108.635 64.420 108.805 64.590 ;
        RECT 108.635 64.060 108.805 64.230 ;
        RECT 110.555 65.620 110.725 65.790 ;
        RECT 110.555 65.260 110.725 65.430 ;
        RECT 110.555 64.900 110.725 65.070 ;
        RECT 110.555 64.540 110.725 64.710 ;
        RECT 110.555 64.180 110.725 64.350 ;
        RECT 111.925 65.620 112.095 65.790 ;
        RECT 111.925 65.260 112.095 65.430 ;
        RECT 111.925 64.900 112.095 65.070 ;
        RECT 111.925 64.540 112.095 64.710 ;
        RECT 111.925 64.180 112.095 64.350 ;
        RECT 113.845 65.670 114.015 65.840 ;
        RECT 113.845 65.310 114.015 65.480 ;
        RECT 113.845 64.950 114.015 65.120 ;
        RECT 113.845 64.590 114.015 64.760 ;
        RECT 113.845 64.230 114.015 64.400 ;
        RECT 108.635 63.700 108.805 63.870 ;
        RECT 109.690 63.760 109.860 63.930 ;
        RECT 110.050 63.760 110.220 63.930 ;
        RECT 111.060 63.760 111.230 63.930 ;
        RECT 111.420 63.760 111.590 63.930 ;
        RECT 112.430 63.760 112.600 63.930 ;
        RECT 112.790 63.760 112.960 63.930 ;
        RECT 113.845 63.870 114.015 64.040 ;
        RECT 113.845 63.510 114.015 63.680 ;
        RECT 108.695 63.090 108.865 63.260 ;
        RECT 109.055 63.090 109.225 63.260 ;
        RECT 109.415 63.090 109.585 63.260 ;
        RECT 109.775 63.090 109.945 63.260 ;
        RECT 110.135 63.090 110.305 63.260 ;
        RECT 110.495 63.090 110.665 63.260 ;
        RECT 110.855 63.090 111.025 63.260 ;
        RECT 111.215 63.090 111.385 63.260 ;
        RECT 111.575 63.090 111.745 63.260 ;
        RECT 111.935 63.090 112.105 63.260 ;
        RECT 112.295 63.090 112.465 63.260 ;
        RECT 112.655 63.090 112.825 63.260 ;
        RECT 113.015 63.090 113.185 63.260 ;
        RECT 113.375 63.090 113.545 63.260 ;
        RECT 113.845 63.150 114.015 63.320 ;
        RECT 114.775 70.570 114.945 70.740 ;
        RECT 115.385 70.630 115.555 70.800 ;
        RECT 115.745 70.630 115.915 70.800 ;
        RECT 116.105 70.630 116.275 70.800 ;
        RECT 116.465 70.630 116.635 70.800 ;
        RECT 116.825 70.630 116.995 70.800 ;
        RECT 117.185 70.630 117.355 70.800 ;
        RECT 114.775 70.210 114.945 70.380 ;
        RECT 114.775 69.850 114.945 70.020 ;
        RECT 115.830 69.960 116.000 70.130 ;
        RECT 116.190 69.960 116.360 70.130 ;
        RECT 117.245 69.950 117.415 70.120 ;
        RECT 114.775 69.490 114.945 69.660 ;
        RECT 114.775 69.130 114.945 69.300 ;
        RECT 114.775 68.770 114.945 68.940 ;
        RECT 114.775 68.410 114.945 68.580 ;
        RECT 114.775 68.050 114.945 68.220 ;
        RECT 116.695 69.540 116.865 69.710 ;
        RECT 116.695 69.180 116.865 69.350 ;
        RECT 116.695 68.820 116.865 68.990 ;
        RECT 116.695 68.460 116.865 68.630 ;
        RECT 116.695 68.100 116.865 68.270 ;
        RECT 117.245 69.590 117.415 69.760 ;
        RECT 117.245 69.230 117.415 69.400 ;
        RECT 117.245 68.870 117.415 69.040 ;
        RECT 117.245 68.510 117.415 68.680 ;
        RECT 117.245 68.150 117.415 68.320 ;
        RECT 114.775 67.690 114.945 67.860 ;
        RECT 115.830 67.680 116.000 67.850 ;
        RECT 116.190 67.680 116.360 67.850 ;
        RECT 117.245 67.790 117.415 67.960 ;
        RECT 114.775 67.330 114.945 67.500 ;
        RECT 117.245 67.430 117.415 67.600 ;
        RECT 114.775 66.970 114.945 67.140 ;
        RECT 114.775 66.610 114.945 66.780 ;
        RECT 114.775 66.250 114.945 66.420 ;
        RECT 114.775 65.890 114.945 66.060 ;
        RECT 115.325 67.260 115.495 67.430 ;
        RECT 115.325 66.900 115.495 67.070 ;
        RECT 115.325 66.540 115.495 66.710 ;
        RECT 115.325 66.180 115.495 66.350 ;
        RECT 115.325 65.820 115.495 65.990 ;
        RECT 117.245 67.070 117.415 67.240 ;
        RECT 117.245 66.710 117.415 66.880 ;
        RECT 117.245 66.350 117.415 66.520 ;
        RECT 117.245 65.990 117.415 66.160 ;
        RECT 117.245 65.630 117.415 65.800 ;
        RECT 115.830 65.400 116.000 65.570 ;
        RECT 116.190 65.400 116.360 65.570 ;
        RECT 118.470 70.290 118.640 70.460 ;
        RECT 119.080 70.350 119.250 70.520 ;
        RECT 119.440 70.350 119.610 70.520 ;
        RECT 119.800 70.350 119.970 70.520 ;
        RECT 120.160 70.350 120.330 70.520 ;
        RECT 120.520 70.350 120.690 70.520 ;
        RECT 120.880 70.350 121.050 70.520 ;
        RECT 121.435 70.350 121.605 70.520 ;
        RECT 121.795 70.350 121.965 70.520 ;
        RECT 122.155 70.350 122.325 70.520 ;
        RECT 122.515 70.350 122.685 70.520 ;
        RECT 122.875 70.350 123.045 70.520 ;
        RECT 123.235 70.350 123.405 70.520 ;
        RECT 123.595 70.350 123.765 70.520 ;
        RECT 118.470 69.930 118.640 70.100 ;
        RECT 123.655 69.950 123.825 70.120 ;
        RECT 118.470 69.570 118.640 69.740 ;
        RECT 119.525 69.680 119.695 69.850 ;
        RECT 119.885 69.680 120.055 69.850 ;
        RECT 122.240 69.680 122.410 69.850 ;
        RECT 122.600 69.680 122.770 69.850 ;
        RECT 123.655 69.590 123.825 69.760 ;
        RECT 118.470 69.210 118.640 69.380 ;
        RECT 119.020 69.250 119.190 69.420 ;
        RECT 119.525 69.250 119.695 69.420 ;
        RECT 119.885 69.250 120.055 69.420 ;
        RECT 121.735 69.250 121.905 69.420 ;
        RECT 122.240 69.250 122.410 69.420 ;
        RECT 122.600 69.250 122.770 69.420 ;
        RECT 118.470 68.850 118.640 69.020 ;
        RECT 123.655 69.230 123.825 69.400 ;
        RECT 119.525 68.820 119.695 68.990 ;
        RECT 119.885 68.820 120.055 68.990 ;
        RECT 122.240 68.820 122.410 68.990 ;
        RECT 122.600 68.820 122.770 68.990 ;
        RECT 123.655 68.870 123.825 69.040 ;
        RECT 118.470 68.490 118.640 68.660 ;
        RECT 119.525 68.390 119.695 68.560 ;
        RECT 119.885 68.390 120.055 68.560 ;
        RECT 120.390 68.390 120.560 68.560 ;
        RECT 122.240 68.390 122.410 68.560 ;
        RECT 122.600 68.390 122.770 68.560 ;
        RECT 123.105 68.390 123.275 68.560 ;
        RECT 123.655 68.510 123.825 68.680 ;
        RECT 118.470 68.130 118.640 68.300 ;
        RECT 123.655 68.150 123.825 68.320 ;
        RECT 119.525 67.960 119.695 68.130 ;
        RECT 119.885 67.960 120.055 68.130 ;
        RECT 122.240 67.960 122.410 68.130 ;
        RECT 122.600 67.960 122.770 68.130 ;
        RECT 118.470 67.770 118.640 67.940 ;
        RECT 123.655 67.790 123.825 67.960 ;
        RECT 118.470 67.410 118.640 67.580 ;
        RECT 119.525 67.530 119.695 67.700 ;
        RECT 119.885 67.530 120.055 67.700 ;
        RECT 120.390 67.530 120.560 67.700 ;
        RECT 122.240 67.530 122.410 67.700 ;
        RECT 122.600 67.530 122.770 67.700 ;
        RECT 123.105 67.530 123.275 67.700 ;
        RECT 123.655 67.430 123.825 67.600 ;
        RECT 118.470 67.050 118.640 67.220 ;
        RECT 119.525 67.100 119.695 67.270 ;
        RECT 119.885 67.100 120.055 67.270 ;
        RECT 122.240 67.100 122.410 67.270 ;
        RECT 122.600 67.100 122.770 67.270 ;
        RECT 118.470 66.690 118.640 66.860 ;
        RECT 123.655 67.070 123.825 67.240 ;
        RECT 119.020 66.670 119.190 66.840 ;
        RECT 119.525 66.670 119.695 66.840 ;
        RECT 119.885 66.670 120.055 66.840 ;
        RECT 121.735 66.670 121.905 66.840 ;
        RECT 122.240 66.670 122.410 66.840 ;
        RECT 122.600 66.670 122.770 66.840 ;
        RECT 123.655 66.710 123.825 66.880 ;
        RECT 118.470 66.330 118.640 66.500 ;
        RECT 119.525 66.240 119.695 66.410 ;
        RECT 119.885 66.240 120.055 66.410 ;
        RECT 122.240 66.240 122.410 66.410 ;
        RECT 122.600 66.240 122.770 66.410 ;
        RECT 123.655 66.350 123.825 66.520 ;
        RECT 118.470 65.970 118.640 66.140 ;
        RECT 123.655 65.990 123.825 66.160 ;
        RECT 118.530 65.570 118.700 65.740 ;
        RECT 118.890 65.570 119.060 65.740 ;
        RECT 119.250 65.570 119.420 65.740 ;
        RECT 119.610 65.570 119.780 65.740 ;
        RECT 119.970 65.570 120.140 65.740 ;
        RECT 120.330 65.570 120.500 65.740 ;
        RECT 120.690 65.570 120.860 65.740 ;
        RECT 121.050 65.570 121.220 65.740 ;
        RECT 121.410 65.570 121.580 65.740 ;
        RECT 121.770 65.570 121.940 65.740 ;
        RECT 122.130 65.570 122.300 65.740 ;
        RECT 122.490 65.570 122.660 65.740 ;
        RECT 122.850 65.570 123.020 65.740 ;
        RECT 123.210 65.570 123.380 65.740 ;
        RECT 123.655 65.630 123.825 65.800 ;
        RECT 124.455 70.250 124.625 70.420 ;
        RECT 125.065 70.310 125.235 70.480 ;
        RECT 125.425 70.310 125.595 70.480 ;
        RECT 125.785 70.310 125.955 70.480 ;
        RECT 126.145 70.310 126.315 70.480 ;
        RECT 126.505 70.310 126.675 70.480 ;
        RECT 126.865 70.310 127.035 70.480 ;
        RECT 124.455 69.890 124.625 70.060 ;
        RECT 126.925 69.870 127.095 70.040 ;
        RECT 124.455 69.530 124.625 69.700 ;
        RECT 125.510 69.680 125.680 69.850 ;
        RECT 125.870 69.680 126.040 69.850 ;
        RECT 126.925 69.510 127.095 69.680 ;
        RECT 124.455 69.170 124.625 69.340 ;
        RECT 125.005 69.250 125.175 69.420 ;
        RECT 125.510 69.250 125.680 69.420 ;
        RECT 125.870 69.250 126.040 69.420 ;
        RECT 126.925 69.150 127.095 69.320 ;
        RECT 124.455 68.810 124.625 68.980 ;
        RECT 125.510 68.820 125.680 68.990 ;
        RECT 125.870 68.820 126.040 68.990 ;
        RECT 124.455 68.450 124.625 68.620 ;
        RECT 126.925 68.790 127.095 68.960 ;
        RECT 125.005 68.390 125.175 68.560 ;
        RECT 125.510 68.390 125.680 68.560 ;
        RECT 125.870 68.390 126.040 68.560 ;
        RECT 126.925 68.430 127.095 68.600 ;
        RECT 124.455 68.090 124.625 68.260 ;
        RECT 125.510 67.960 125.680 68.130 ;
        RECT 125.870 67.960 126.040 68.130 ;
        RECT 126.925 68.070 127.095 68.240 ;
        RECT 124.455 67.730 124.625 67.900 ;
        RECT 126.925 67.710 127.095 67.880 ;
        RECT 124.455 67.370 124.625 67.540 ;
        RECT 125.005 67.530 125.175 67.700 ;
        RECT 125.510 67.530 125.680 67.700 ;
        RECT 125.870 67.530 126.040 67.700 ;
        RECT 126.925 67.350 127.095 67.520 ;
        RECT 124.455 67.010 124.625 67.180 ;
        RECT 125.510 67.100 125.680 67.270 ;
        RECT 125.870 67.100 126.040 67.270 ;
        RECT 126.925 66.990 127.095 67.160 ;
        RECT 124.455 66.650 124.625 66.820 ;
        RECT 125.005 66.670 125.175 66.840 ;
        RECT 125.510 66.670 125.680 66.840 ;
        RECT 125.870 66.670 126.040 66.840 ;
        RECT 124.455 66.290 124.625 66.460 ;
        RECT 126.925 66.630 127.095 66.800 ;
        RECT 125.510 66.240 125.680 66.410 ;
        RECT 125.870 66.240 126.040 66.410 ;
        RECT 126.925 66.270 127.095 66.440 ;
        RECT 124.455 65.930 124.625 66.100 ;
        RECT 125.510 65.810 125.680 65.980 ;
        RECT 125.870 65.810 126.040 65.980 ;
        RECT 126.375 65.810 126.545 65.980 ;
        RECT 126.925 65.910 127.095 66.080 ;
        RECT 124.455 65.570 124.625 65.740 ;
        RECT 114.775 65.220 114.945 65.390 ;
        RECT 117.245 65.270 117.415 65.440 ;
        RECT 114.775 64.860 114.945 65.030 ;
        RECT 114.775 64.500 114.945 64.670 ;
        RECT 114.775 64.140 114.945 64.310 ;
        RECT 114.775 63.780 114.945 63.950 ;
        RECT 114.775 63.420 114.945 63.590 ;
        RECT 115.325 64.980 115.495 65.150 ;
        RECT 115.325 64.620 115.495 64.790 ;
        RECT 115.325 64.260 115.495 64.430 ;
        RECT 115.325 63.900 115.495 64.070 ;
        RECT 115.325 63.540 115.495 63.710 ;
        RECT 126.925 65.550 127.095 65.720 ;
        RECT 125.510 65.380 125.680 65.550 ;
        RECT 125.870 65.380 126.040 65.550 ;
        RECT 117.245 64.910 117.415 65.080 ;
        RECT 117.245 64.550 117.415 64.720 ;
        RECT 117.245 64.190 117.415 64.360 ;
        RECT 117.245 63.830 117.415 64.000 ;
        RECT 117.245 63.470 117.415 63.640 ;
        RECT 114.775 63.060 114.945 63.230 ;
        RECT 115.830 63.120 116.000 63.290 ;
        RECT 116.190 63.120 116.360 63.290 ;
        RECT 117.245 63.110 117.415 63.280 ;
        RECT 114.775 62.700 114.945 62.870 ;
        RECT 114.775 62.340 114.945 62.510 ;
        RECT 114.775 61.980 114.945 62.150 ;
        RECT 114.775 61.620 114.945 61.790 ;
        RECT 114.775 61.260 114.945 61.430 ;
        RECT 116.695 62.700 116.865 62.870 ;
        RECT 116.695 62.340 116.865 62.510 ;
        RECT 116.695 61.980 116.865 62.150 ;
        RECT 116.695 61.620 116.865 61.790 ;
        RECT 116.695 61.260 116.865 61.430 ;
        RECT 117.245 62.750 117.415 62.920 ;
        RECT 117.245 62.390 117.415 62.560 ;
        RECT 117.245 62.030 117.415 62.200 ;
        RECT 117.245 61.670 117.415 61.840 ;
        RECT 117.245 61.310 117.415 61.480 ;
        RECT 114.775 60.900 114.945 61.070 ;
        RECT 115.830 60.840 116.000 61.010 ;
        RECT 116.190 60.840 116.360 61.010 ;
        RECT 117.245 60.950 117.415 61.120 ;
        RECT 114.775 60.540 114.945 60.710 ;
        RECT 117.245 60.590 117.415 60.760 ;
        RECT 114.835 60.170 115.005 60.340 ;
        RECT 115.195 60.170 115.365 60.340 ;
        RECT 115.555 60.170 115.725 60.340 ;
        RECT 115.915 60.170 116.085 60.340 ;
        RECT 116.275 60.170 116.445 60.340 ;
        RECT 116.635 60.170 116.805 60.340 ;
        RECT 117.245 60.230 117.415 60.400 ;
        RECT 118.470 65.000 118.640 65.170 ;
        RECT 119.080 65.060 119.250 65.230 ;
        RECT 119.440 65.060 119.610 65.230 ;
        RECT 119.800 65.060 119.970 65.230 ;
        RECT 120.160 65.060 120.330 65.230 ;
        RECT 120.520 65.060 120.690 65.230 ;
        RECT 120.880 65.060 121.050 65.230 ;
        RECT 121.435 65.060 121.605 65.230 ;
        RECT 121.795 65.060 121.965 65.230 ;
        RECT 122.155 65.060 122.325 65.230 ;
        RECT 122.515 65.060 122.685 65.230 ;
        RECT 122.875 65.060 123.045 65.230 ;
        RECT 123.235 65.060 123.405 65.230 ;
        RECT 123.595 65.060 123.765 65.230 ;
        RECT 118.470 64.640 118.640 64.810 ;
        RECT 118.470 64.280 118.640 64.450 ;
        RECT 119.525 64.430 119.695 64.600 ;
        RECT 119.885 64.430 120.055 64.600 ;
        RECT 122.240 64.430 122.410 64.600 ;
        RECT 122.600 64.430 122.770 64.600 ;
        RECT 123.655 64.380 123.825 64.550 ;
        RECT 118.470 63.920 118.640 64.090 ;
        RECT 119.020 64.000 119.190 64.170 ;
        RECT 119.525 64.000 119.695 64.170 ;
        RECT 119.885 64.000 120.055 64.170 ;
        RECT 121.735 64.000 121.905 64.170 ;
        RECT 122.240 64.000 122.410 64.170 ;
        RECT 122.600 64.000 122.770 64.170 ;
        RECT 123.655 64.020 123.825 64.190 ;
        RECT 118.470 63.560 118.640 63.730 ;
        RECT 119.525 63.570 119.695 63.740 ;
        RECT 119.885 63.570 120.055 63.740 ;
        RECT 122.240 63.570 122.410 63.740 ;
        RECT 122.600 63.570 122.770 63.740 ;
        RECT 123.655 63.660 123.825 63.830 ;
        RECT 118.470 63.200 118.640 63.370 ;
        RECT 119.525 63.140 119.695 63.310 ;
        RECT 119.885 63.140 120.055 63.310 ;
        RECT 120.390 63.140 120.560 63.310 ;
        RECT 122.240 63.140 122.410 63.310 ;
        RECT 122.600 63.140 122.770 63.310 ;
        RECT 123.105 63.140 123.275 63.310 ;
        RECT 123.655 63.300 123.825 63.470 ;
        RECT 118.470 62.840 118.640 63.010 ;
        RECT 123.655 62.940 123.825 63.110 ;
        RECT 119.525 62.710 119.695 62.880 ;
        RECT 119.885 62.710 120.055 62.880 ;
        RECT 122.240 62.710 122.410 62.880 ;
        RECT 122.600 62.710 122.770 62.880 ;
        RECT 118.470 62.480 118.640 62.650 ;
        RECT 123.655 62.580 123.825 62.750 ;
        RECT 118.470 62.120 118.640 62.290 ;
        RECT 119.525 62.280 119.695 62.450 ;
        RECT 119.885 62.280 120.055 62.450 ;
        RECT 120.390 62.280 120.560 62.450 ;
        RECT 122.240 62.280 122.410 62.450 ;
        RECT 122.600 62.280 122.770 62.450 ;
        RECT 123.105 62.280 123.275 62.450 ;
        RECT 123.655 62.220 123.825 62.390 ;
        RECT 118.470 61.760 118.640 61.930 ;
        RECT 119.525 61.850 119.695 62.020 ;
        RECT 119.885 61.850 120.055 62.020 ;
        RECT 122.240 61.850 122.410 62.020 ;
        RECT 122.600 61.850 122.770 62.020 ;
        RECT 123.655 61.860 123.825 62.030 ;
        RECT 118.470 61.400 118.640 61.570 ;
        RECT 119.020 61.420 119.190 61.590 ;
        RECT 119.525 61.420 119.695 61.590 ;
        RECT 119.885 61.420 120.055 61.590 ;
        RECT 121.735 61.420 121.905 61.590 ;
        RECT 122.240 61.420 122.410 61.590 ;
        RECT 122.600 61.420 122.770 61.590 ;
        RECT 123.655 61.500 123.825 61.670 ;
        RECT 118.470 61.040 118.640 61.210 ;
        RECT 119.525 60.990 119.695 61.160 ;
        RECT 119.885 60.990 120.055 61.160 ;
        RECT 122.240 60.990 122.410 61.160 ;
        RECT 122.600 60.990 122.770 61.160 ;
        RECT 123.655 61.140 123.825 61.310 ;
        RECT 123.655 60.780 123.825 60.950 ;
        RECT 118.530 60.360 118.700 60.530 ;
        RECT 118.890 60.360 119.060 60.530 ;
        RECT 119.250 60.360 119.420 60.530 ;
        RECT 119.610 60.360 119.780 60.530 ;
        RECT 119.970 60.360 120.140 60.530 ;
        RECT 120.330 60.360 120.500 60.530 ;
        RECT 120.690 60.360 120.860 60.530 ;
        RECT 121.050 60.360 121.220 60.530 ;
        RECT 121.410 60.360 121.580 60.530 ;
        RECT 121.770 60.360 121.940 60.530 ;
        RECT 122.130 60.360 122.300 60.530 ;
        RECT 122.490 60.360 122.660 60.530 ;
        RECT 122.850 60.360 123.020 60.530 ;
        RECT 123.210 60.360 123.380 60.530 ;
        RECT 123.655 60.420 123.825 60.590 ;
        RECT 124.455 65.200 124.625 65.370 ;
        RECT 126.925 65.190 127.095 65.360 ;
        RECT 124.455 64.840 124.625 65.010 ;
        RECT 125.510 64.950 125.680 65.120 ;
        RECT 125.870 64.950 126.040 65.120 ;
        RECT 126.375 64.950 126.545 65.120 ;
        RECT 126.925 64.830 127.095 65.000 ;
        RECT 124.455 64.480 124.625 64.650 ;
        RECT 125.510 64.520 125.680 64.690 ;
        RECT 125.870 64.520 126.040 64.690 ;
        RECT 124.455 64.120 124.625 64.290 ;
        RECT 126.925 64.470 127.095 64.640 ;
        RECT 125.005 64.090 125.175 64.260 ;
        RECT 125.510 64.090 125.680 64.260 ;
        RECT 125.870 64.090 126.040 64.260 ;
        RECT 126.925 64.110 127.095 64.280 ;
        RECT 124.455 63.760 124.625 63.930 ;
        RECT 125.510 63.660 125.680 63.830 ;
        RECT 125.870 63.660 126.040 63.830 ;
        RECT 126.925 63.750 127.095 63.920 ;
        RECT 124.455 63.400 124.625 63.570 ;
        RECT 125.005 63.230 125.175 63.400 ;
        RECT 125.510 63.230 125.680 63.400 ;
        RECT 125.870 63.230 126.040 63.400 ;
        RECT 126.925 63.390 127.095 63.560 ;
        RECT 124.455 63.040 124.625 63.210 ;
        RECT 126.925 63.030 127.095 63.200 ;
        RECT 124.455 62.680 124.625 62.850 ;
        RECT 125.510 62.800 125.680 62.970 ;
        RECT 125.870 62.800 126.040 62.970 ;
        RECT 126.925 62.670 127.095 62.840 ;
        RECT 124.455 62.320 124.625 62.490 ;
        RECT 125.005 62.370 125.175 62.540 ;
        RECT 125.510 62.370 125.680 62.540 ;
        RECT 125.870 62.370 126.040 62.540 ;
        RECT 124.455 61.960 124.625 62.130 ;
        RECT 126.925 62.310 127.095 62.480 ;
        RECT 125.510 61.940 125.680 62.110 ;
        RECT 125.870 61.940 126.040 62.110 ;
        RECT 126.925 61.950 127.095 62.120 ;
        RECT 124.455 61.600 124.625 61.770 ;
        RECT 125.005 61.510 125.175 61.680 ;
        RECT 125.510 61.510 125.680 61.680 ;
        RECT 125.870 61.510 126.040 61.680 ;
        RECT 126.925 61.590 127.095 61.760 ;
        RECT 124.455 61.240 124.625 61.410 ;
        RECT 125.510 61.080 125.680 61.250 ;
        RECT 125.870 61.080 126.040 61.250 ;
        RECT 126.925 61.230 127.095 61.400 ;
        RECT 124.455 60.880 124.625 61.050 ;
        RECT 126.925 60.870 127.095 61.040 ;
        RECT 124.515 60.450 124.685 60.620 ;
        RECT 124.875 60.450 125.045 60.620 ;
        RECT 125.235 60.450 125.405 60.620 ;
        RECT 125.595 60.450 125.765 60.620 ;
        RECT 125.955 60.450 126.125 60.620 ;
        RECT 126.315 60.450 126.485 60.620 ;
        RECT 126.925 60.510 127.095 60.680 ;
      LAYER met1 ;
        RECT 107.530 173.840 110.225 174.130 ;
        RECT 110.515 173.840 114.235 174.130 ;
        RECT 107.530 169.350 107.820 173.840 ;
        RECT 108.195 173.185 109.195 173.445 ;
        RECT 108.195 172.755 109.195 173.015 ;
        RECT 109.385 172.590 109.675 173.840 ;
        RECT 108.195 172.325 109.195 172.585 ;
        RECT 108.195 171.895 109.195 172.155 ;
        RECT 109.385 171.760 109.675 172.320 ;
        RECT 110.205 171.760 110.535 173.435 ;
        RECT 111.065 172.590 111.355 173.840 ;
        RECT 112.045 173.430 113.045 173.445 ;
        RECT 111.545 173.200 113.545 173.430 ;
        RECT 112.045 173.185 113.045 173.200 ;
        RECT 112.045 173.000 113.045 173.015 ;
        RECT 111.545 172.770 113.545 173.000 ;
        RECT 112.045 172.755 113.045 172.770 ;
        RECT 112.045 172.570 113.045 172.585 ;
        RECT 111.545 172.340 113.545 172.570 ;
        RECT 112.045 172.325 113.045 172.340 ;
        RECT 111.065 171.760 111.355 172.320 ;
        RECT 111.545 171.895 113.545 172.155 ;
        RECT 108.195 171.465 109.195 171.725 ;
        RECT 109.385 171.430 111.355 171.760 ;
        RECT 112.045 171.710 113.045 171.725 ;
        RECT 111.545 171.480 113.545 171.710 ;
        RECT 112.045 171.465 113.045 171.480 ;
        RECT 108.195 171.035 109.195 171.295 ;
        RECT 109.385 170.870 109.675 171.430 ;
        RECT 111.065 170.870 111.355 171.430 ;
        RECT 111.545 171.035 113.545 171.295 ;
        RECT 108.195 170.605 109.195 170.865 ;
        RECT 112.045 170.850 113.045 170.865 ;
        RECT 111.545 170.620 113.545 170.850 ;
        RECT 112.045 170.605 113.045 170.620 ;
        RECT 108.195 170.175 109.195 170.435 ;
        RECT 108.195 169.745 109.195 170.005 ;
        RECT 109.385 169.350 109.675 170.600 ;
        RECT 111.065 169.350 111.355 170.600 ;
        RECT 112.045 170.420 113.045 170.435 ;
        RECT 111.545 170.190 113.545 170.420 ;
        RECT 112.045 170.175 113.045 170.190 ;
        RECT 112.045 169.990 113.045 170.005 ;
        RECT 111.545 169.760 113.545 169.990 ;
        RECT 112.045 169.745 113.045 169.760 ;
        RECT 113.945 169.350 114.235 173.840 ;
        RECT 107.530 169.060 110.225 169.350 ;
        RECT 110.515 169.060 114.235 169.350 ;
        RECT 108.575 164.690 114.075 164.980 ;
        RECT 56.120 151.440 62.770 151.730 ;
        RECT 56.120 112.230 56.410 151.440 ;
        RECT 57.150 141.545 58.150 141.805 ;
        RECT 57.150 139.265 58.150 139.525 ;
        RECT 57.150 136.985 58.150 137.245 ;
        RECT 57.150 134.705 58.150 134.965 ;
        RECT 57.150 132.425 58.150 132.685 ;
        RECT 58.340 130.580 58.630 151.440 ;
        RECT 60.260 149.660 60.550 151.440 ;
        RECT 60.740 150.785 61.740 151.045 ;
        RECT 60.740 150.005 61.740 150.265 ;
        RECT 60.740 149.225 61.740 149.485 ;
        RECT 60.740 146.945 61.740 147.205 ;
        RECT 61.930 145.100 62.260 149.050 ;
        RECT 60.740 144.665 61.740 144.925 ;
        RECT 60.260 144.160 60.550 144.490 ;
        RECT 60.260 143.870 61.740 144.160 ;
        RECT 60.260 143.380 60.550 143.870 ;
        RECT 60.260 143.090 61.740 143.380 ;
        RECT 60.260 142.600 60.550 143.090 ;
        RECT 60.260 142.310 61.740 142.600 ;
        RECT 60.260 141.980 60.550 142.310 ;
        RECT 60.740 141.545 61.740 141.805 ;
        RECT 60.260 139.700 60.550 141.370 ;
        RECT 60.740 139.265 61.740 139.525 ;
        RECT 60.260 137.420 60.550 139.090 ;
        RECT 60.740 136.985 61.740 137.245 ;
        RECT 60.260 135.140 60.550 136.810 ;
        RECT 60.740 134.705 61.740 134.965 ;
        RECT 60.260 132.860 60.550 134.530 ;
        RECT 60.740 132.425 61.740 132.685 ;
        RECT 60.260 130.580 60.550 132.250 ;
        RECT 57.150 130.145 58.150 130.405 ;
        RECT 60.740 130.145 61.740 130.405 ;
        RECT 56.630 126.020 56.960 129.970 ;
        RECT 60.260 128.300 60.550 129.970 ;
        RECT 61.930 128.300 62.260 141.370 ;
        RECT 57.150 127.865 58.150 128.125 ;
        RECT 60.740 127.865 61.740 128.125 ;
        RECT 60.260 126.020 60.550 127.690 ;
        RECT 57.150 125.585 58.150 125.845 ;
        RECT 60.740 125.585 61.740 125.845 ;
        RECT 57.150 123.305 58.150 123.565 ;
        RECT 57.150 121.025 58.150 121.285 ;
        RECT 57.150 118.745 58.150 119.005 ;
        RECT 57.150 116.465 58.150 116.725 ;
        RECT 57.150 114.185 58.150 114.445 ;
        RECT 58.340 112.230 58.630 125.410 ;
        RECT 60.260 123.740 60.550 125.410 ;
        RECT 60.740 123.305 61.740 123.565 ;
        RECT 60.260 121.460 60.550 123.130 ;
        RECT 60.740 121.025 61.740 121.285 ;
        RECT 60.260 119.180 60.550 120.850 ;
        RECT 60.740 118.745 61.740 119.005 ;
        RECT 60.260 116.900 60.550 118.570 ;
        RECT 60.740 116.465 61.740 116.725 ;
        RECT 60.260 114.620 60.550 116.290 ;
        RECT 61.930 114.620 62.260 127.690 ;
        RECT 60.740 114.185 61.740 114.445 ;
        RECT 60.260 112.230 60.550 114.010 ;
        RECT 60.740 113.405 61.740 113.665 ;
        RECT 60.740 112.625 61.740 112.885 ;
        RECT 62.480 112.230 62.770 151.440 ;
        RECT 64.375 151.440 66.935 151.730 ;
        RECT 64.375 142.710 64.665 151.440 ;
        RECT 65.405 150.785 65.905 151.045 ;
        RECT 65.405 150.005 65.905 150.265 ;
        RECT 66.095 149.660 66.385 151.440 ;
        RECT 65.405 149.225 65.905 149.485 ;
        RECT 64.885 145.100 65.215 149.050 ;
        RECT 65.405 146.945 65.905 147.205 ;
        RECT 65.405 144.665 65.905 144.925 ;
        RECT 65.405 143.885 65.905 144.145 ;
        RECT 65.405 143.105 65.905 143.365 ;
        RECT 66.095 142.710 66.385 144.490 ;
        RECT 66.645 142.710 66.935 151.440 ;
        RECT 91.855 151.440 94.415 151.730 ;
        RECT 64.375 142.420 66.935 142.710 ;
        RECT 72.530 142.720 77.830 143.010 ;
        RECT 64.375 138.230 66.935 138.520 ;
        RECT 64.375 117.820 64.665 138.230 ;
        RECT 64.925 135.405 65.215 138.230 ;
        RECT 65.405 137.575 65.905 137.835 ;
        RECT 66.075 137.435 66.365 138.230 ;
        RECT 65.405 136.295 65.905 136.555 ;
        RECT 66.075 135.405 66.385 137.435 ;
        RECT 65.405 135.015 65.905 135.275 ;
        RECT 64.885 133.015 65.215 134.975 ;
        RECT 66.095 133.015 66.425 134.840 ;
        RECT 64.885 132.725 66.425 133.015 ;
        RECT 64.885 130.890 65.215 132.725 ;
        RECT 66.095 130.890 66.425 132.725 ;
        RECT 65.405 130.455 65.905 130.715 ;
        RECT 64.925 129.445 65.215 130.315 ;
        RECT 66.075 129.445 66.385 130.315 ;
        RECT 64.925 129.165 66.385 129.445 ;
        RECT 64.925 128.165 65.215 129.165 ;
        RECT 66.075 128.285 66.385 129.165 ;
        RECT 66.075 128.165 66.365 128.285 ;
        RECT 64.925 127.885 66.365 128.165 ;
        RECT 64.925 126.885 65.215 127.885 ;
        RECT 66.075 127.755 66.365 127.885 ;
        RECT 66.075 126.885 66.385 127.755 ;
        RECT 64.925 126.605 66.385 126.885 ;
        RECT 64.925 125.725 65.215 126.605 ;
        RECT 66.075 125.725 66.385 126.605 ;
        RECT 65.405 125.335 65.905 125.595 ;
        RECT 64.880 123.490 65.215 125.160 ;
        RECT 64.880 122.880 65.210 123.490 ;
        RECT 65.405 123.055 65.905 123.315 ;
        RECT 64.880 121.210 65.215 122.880 ;
        RECT 65.405 120.775 65.905 121.035 ;
        RECT 64.925 117.820 65.215 120.635 ;
        RECT 65.405 119.495 65.905 119.755 ;
        RECT 66.075 118.605 66.385 120.635 ;
        RECT 65.405 118.215 65.905 118.475 ;
        RECT 66.075 117.820 66.365 118.605 ;
        RECT 66.645 117.820 66.935 138.230 ;
        RECT 64.375 117.530 66.935 117.820 ;
        RECT 68.130 138.230 71.190 138.520 ;
        RECT 68.130 117.820 68.420 138.230 ;
        RECT 68.700 137.435 68.990 138.230 ;
        RECT 69.160 137.575 70.160 137.835 ;
        RECT 68.680 135.405 68.990 137.435 ;
        RECT 70.330 137.435 70.620 138.230 ;
        RECT 69.160 136.295 70.160 136.555 ;
        RECT 70.330 135.405 70.640 137.435 ;
        RECT 69.160 135.015 70.160 135.275 ;
        RECT 68.640 130.890 68.970 134.840 ;
        RECT 70.330 132.980 70.660 134.840 ;
        RECT 69.160 132.715 70.660 132.980 ;
        RECT 70.330 130.890 70.660 132.715 ;
        RECT 69.160 130.455 70.160 130.715 ;
        RECT 68.680 129.445 68.990 130.315 ;
        RECT 70.330 129.445 70.640 130.315 ;
        RECT 68.680 129.165 70.640 129.445 ;
        RECT 68.680 128.285 68.990 129.165 ;
        RECT 68.700 128.165 68.990 128.285 ;
        RECT 70.330 128.285 70.640 129.165 ;
        RECT 70.330 128.165 70.620 128.285 ;
        RECT 68.700 127.885 70.620 128.165 ;
        RECT 68.700 127.755 68.990 127.885 ;
        RECT 68.680 126.885 68.990 127.755 ;
        RECT 70.330 127.755 70.620 127.885 ;
        RECT 70.330 126.885 70.640 127.755 ;
        RECT 68.680 126.605 70.640 126.885 ;
        RECT 68.680 125.725 68.990 126.605 ;
        RECT 70.330 125.725 70.640 126.605 ;
        RECT 69.160 125.335 70.160 125.595 ;
        RECT 70.330 123.300 70.660 125.160 ;
        RECT 69.160 123.025 70.660 123.300 ;
        RECT 70.330 121.210 70.660 123.025 ;
        RECT 69.160 120.775 70.160 121.035 ;
        RECT 68.680 118.605 68.990 120.635 ;
        RECT 69.160 119.495 70.160 119.755 ;
        RECT 68.700 117.820 68.990 118.605 ;
        RECT 70.330 118.605 70.640 120.635 ;
        RECT 69.160 118.215 70.160 118.475 ;
        RECT 70.330 117.820 70.620 118.605 ;
        RECT 70.900 117.820 71.190 138.230 ;
        RECT 68.130 117.530 71.190 117.820 ;
        RECT 56.120 111.940 62.770 112.230 ;
        RECT 63.625 113.280 67.345 113.570 ;
        RECT 67.610 113.280 70.305 113.570 ;
        RECT 63.625 89.430 63.915 113.280 ;
        RECT 64.315 112.625 65.315 112.885 ;
        RECT 64.315 110.345 65.315 110.605 ;
        RECT 65.505 108.500 65.795 113.280 ;
        RECT 68.635 108.500 68.925 113.280 ;
        RECT 69.115 112.625 69.615 112.885 ;
        RECT 69.115 110.345 69.615 110.605 ;
        RECT 64.315 108.065 65.315 108.325 ;
        RECT 69.115 108.065 69.615 108.325 ;
        RECT 64.315 105.785 65.315 106.045 ;
        RECT 65.505 103.940 65.835 107.890 ;
        RECT 67.025 105.775 67.985 106.055 ;
        RECT 64.315 103.505 65.315 103.765 ;
        RECT 67.340 103.330 67.670 105.775 ;
        RECT 68.595 103.940 68.925 107.890 ;
        RECT 69.115 105.785 69.615 106.045 ;
        RECT 69.115 103.505 69.615 103.765 ;
        RECT 65.505 103.000 68.925 103.330 ;
        RECT 64.315 101.225 65.315 101.485 ;
        RECT 65.505 99.380 65.835 103.000 ;
        RECT 67.025 101.215 67.985 101.495 ;
        RECT 64.315 98.945 65.315 99.205 ;
        RECT 67.340 98.770 67.670 101.215 ;
        RECT 68.595 99.380 68.925 103.000 ;
        RECT 69.115 101.225 69.615 101.485 ;
        RECT 69.115 98.945 69.615 99.205 ;
        RECT 65.505 98.440 68.925 98.770 ;
        RECT 64.315 96.665 65.315 96.925 ;
        RECT 65.505 94.820 65.835 98.440 ;
        RECT 68.595 94.820 68.925 98.440 ;
        RECT 69.115 96.665 69.615 96.925 ;
        RECT 64.315 94.385 65.315 94.645 ;
        RECT 69.115 94.385 69.615 94.645 ;
        RECT 64.315 92.105 65.315 92.365 ;
        RECT 64.315 89.825 65.315 90.085 ;
        RECT 65.505 89.430 65.795 94.210 ;
        RECT 68.635 89.430 68.925 94.210 ;
        RECT 69.115 92.105 69.615 92.365 ;
        RECT 69.115 89.825 69.615 90.085 ;
        RECT 70.015 89.430 70.305 113.280 ;
        RECT 72.530 113.270 72.820 142.720 ;
        RECT 73.560 142.105 74.060 142.365 ;
        RECT 73.040 130.860 73.370 141.370 ;
        RECT 74.250 141.070 74.540 142.720 ;
        RECT 73.560 140.840 74.540 141.070 ;
        RECT 74.250 139.935 74.540 140.840 ;
        RECT 73.560 139.545 74.060 139.805 ;
        RECT 74.250 137.700 74.540 139.370 ;
        RECT 73.560 137.265 74.060 137.525 ;
        RECT 74.250 135.420 74.540 137.090 ;
        RECT 75.820 135.535 76.110 142.720 ;
        RECT 76.300 141.705 76.800 141.965 ;
        RECT 76.300 138.425 76.800 138.685 ;
        RECT 76.990 135.535 77.280 142.720 ;
        RECT 73.560 134.985 74.060 135.245 ;
        RECT 76.300 135.145 76.800 135.405 ;
        RECT 74.250 133.140 74.540 134.810 ;
        RECT 73.560 132.705 74.060 132.965 ;
        RECT 74.250 130.860 74.540 132.530 ;
        RECT 73.560 130.425 74.060 130.685 ;
        RECT 73.080 129.415 73.370 130.285 ;
        RECT 74.250 129.415 74.540 130.285 ;
        RECT 73.080 129.135 74.540 129.415 ;
        RECT 73.080 128.135 73.370 129.135 ;
        RECT 74.250 128.135 74.540 129.135 ;
        RECT 73.080 127.855 74.540 128.135 ;
        RECT 76.300 127.865 76.800 128.125 ;
        RECT 73.080 126.855 73.370 127.855 ;
        RECT 74.250 126.855 74.540 127.855 ;
        RECT 73.080 126.575 74.540 126.855 ;
        RECT 73.080 125.695 73.370 126.575 ;
        RECT 74.250 125.695 74.540 126.575 ;
        RECT 73.560 125.305 74.060 125.565 ;
        RECT 73.040 114.620 73.370 125.130 ;
        RECT 74.250 123.460 74.540 125.130 ;
        RECT 73.560 123.025 74.060 123.285 ;
        RECT 74.250 121.180 74.540 122.850 ;
        RECT 73.560 120.745 74.060 121.005 ;
        RECT 76.990 121.000 77.320 134.990 ;
        RECT 76.300 120.585 76.800 120.845 ;
        RECT 74.250 118.900 74.540 120.570 ;
        RECT 73.560 118.465 74.060 118.725 ;
        RECT 74.250 116.620 74.540 118.290 ;
        RECT 73.560 116.185 74.060 116.445 ;
        RECT 74.250 115.150 74.540 116.045 ;
        RECT 73.560 114.920 74.540 115.150 ;
        RECT 73.560 113.625 74.060 113.885 ;
        RECT 74.250 113.270 74.540 114.920 ;
        RECT 75.820 113.270 76.110 120.445 ;
        RECT 76.300 117.305 76.800 117.565 ;
        RECT 76.300 114.025 76.800 114.285 ;
        RECT 76.990 113.270 77.280 120.445 ;
        RECT 77.540 113.270 77.830 142.720 ;
        RECT 72.530 112.980 77.830 113.270 ;
        RECT 80.960 142.720 86.260 143.010 ;
        RECT 80.960 113.270 81.250 142.720 ;
        RECT 81.510 135.535 81.800 142.720 ;
        RECT 81.990 141.705 82.490 141.965 ;
        RECT 81.990 138.425 82.490 138.685 ;
        RECT 82.680 135.535 82.970 142.720 ;
        RECT 84.250 141.070 84.540 142.720 ;
        RECT 84.730 142.105 85.230 142.365 ;
        RECT 84.250 140.840 85.230 141.070 ;
        RECT 84.250 139.935 84.540 140.840 ;
        RECT 84.730 139.545 85.230 139.805 ;
        RECT 84.250 137.700 84.540 139.370 ;
        RECT 84.730 137.265 85.230 137.525 ;
        RECT 84.250 135.420 84.540 137.090 ;
        RECT 81.990 135.145 82.490 135.405 ;
        RECT 81.470 121.000 81.800 134.990 ;
        RECT 84.730 134.985 85.230 135.245 ;
        RECT 84.250 133.140 84.540 134.810 ;
        RECT 84.730 132.705 85.230 132.965 ;
        RECT 84.250 130.860 84.540 132.530 ;
        RECT 85.420 130.860 85.750 141.370 ;
        RECT 84.730 130.425 85.230 130.685 ;
        RECT 84.250 129.415 84.540 130.285 ;
        RECT 85.420 129.415 85.710 130.285 ;
        RECT 84.250 129.135 85.710 129.415 ;
        RECT 84.250 128.135 84.540 129.135 ;
        RECT 85.420 128.135 85.710 129.135 ;
        RECT 81.990 127.865 82.490 128.125 ;
        RECT 84.250 127.855 85.710 128.135 ;
        RECT 84.250 126.855 84.540 127.855 ;
        RECT 85.420 126.855 85.710 127.855 ;
        RECT 84.250 126.575 85.710 126.855 ;
        RECT 84.250 125.695 84.540 126.575 ;
        RECT 85.420 125.695 85.710 126.575 ;
        RECT 84.730 125.305 85.230 125.565 ;
        RECT 84.250 123.460 84.540 125.130 ;
        RECT 84.730 123.025 85.230 123.285 ;
        RECT 84.250 121.180 84.540 122.850 ;
        RECT 81.990 120.585 82.490 120.845 ;
        RECT 84.730 120.745 85.230 121.005 ;
        RECT 81.510 113.270 81.800 120.445 ;
        RECT 81.990 117.305 82.490 117.565 ;
        RECT 81.990 114.025 82.490 114.285 ;
        RECT 82.680 113.270 82.970 120.445 ;
        RECT 84.250 118.900 84.540 120.570 ;
        RECT 84.730 118.465 85.230 118.725 ;
        RECT 84.250 116.620 84.540 118.290 ;
        RECT 84.730 116.185 85.230 116.445 ;
        RECT 84.250 115.150 84.540 116.045 ;
        RECT 84.250 114.920 85.230 115.150 ;
        RECT 84.250 113.270 84.540 114.920 ;
        RECT 85.420 114.620 85.750 125.130 ;
        RECT 84.730 113.625 85.230 113.885 ;
        RECT 85.970 113.270 86.260 142.720 ;
        RECT 91.855 142.710 92.145 151.440 ;
        RECT 92.405 149.660 92.695 151.440 ;
        RECT 92.885 150.785 93.385 151.045 ;
        RECT 92.885 150.005 93.385 150.265 ;
        RECT 92.885 149.225 93.385 149.485 ;
        RECT 92.885 146.945 93.385 147.205 ;
        RECT 93.575 145.100 93.905 149.050 ;
        RECT 92.885 144.665 93.385 144.925 ;
        RECT 92.405 142.710 92.695 144.490 ;
        RECT 92.885 143.885 93.385 144.145 ;
        RECT 92.885 143.105 93.385 143.365 ;
        RECT 94.125 142.710 94.415 151.440 ;
        RECT 91.855 142.420 94.415 142.710 ;
        RECT 96.020 151.440 102.670 151.730 ;
        RECT 87.600 138.230 90.660 138.520 ;
        RECT 87.600 117.820 87.890 138.230 ;
        RECT 88.170 137.435 88.460 138.230 ;
        RECT 88.630 137.575 89.630 137.835 ;
        RECT 88.150 135.405 88.460 137.435 ;
        RECT 89.800 137.435 90.090 138.230 ;
        RECT 88.630 136.295 89.630 136.555 ;
        RECT 89.800 135.405 90.110 137.435 ;
        RECT 88.630 135.015 89.630 135.275 ;
        RECT 88.130 132.980 88.460 134.840 ;
        RECT 88.130 132.715 89.630 132.980 ;
        RECT 88.130 130.890 88.460 132.715 ;
        RECT 89.820 130.890 90.150 134.840 ;
        RECT 88.630 130.455 89.630 130.715 ;
        RECT 88.150 129.445 88.460 130.315 ;
        RECT 89.800 129.445 90.110 130.315 ;
        RECT 88.150 129.165 90.110 129.445 ;
        RECT 88.150 128.285 88.460 129.165 ;
        RECT 88.170 128.165 88.460 128.285 ;
        RECT 89.800 128.285 90.110 129.165 ;
        RECT 89.800 128.165 90.090 128.285 ;
        RECT 88.170 127.885 90.090 128.165 ;
        RECT 88.170 127.755 88.460 127.885 ;
        RECT 88.150 126.885 88.460 127.755 ;
        RECT 89.800 127.755 90.090 127.885 ;
        RECT 89.800 126.885 90.110 127.755 ;
        RECT 88.150 126.605 90.110 126.885 ;
        RECT 88.150 125.725 88.460 126.605 ;
        RECT 89.800 125.725 90.110 126.605 ;
        RECT 88.630 125.335 89.630 125.595 ;
        RECT 88.130 123.300 88.460 125.160 ;
        RECT 88.130 123.025 89.630 123.300 ;
        RECT 88.130 121.210 88.460 123.025 ;
        RECT 88.630 120.775 89.630 121.035 ;
        RECT 88.150 118.605 88.460 120.635 ;
        RECT 88.630 119.495 89.630 119.755 ;
        RECT 88.170 117.820 88.460 118.605 ;
        RECT 89.800 118.605 90.110 120.635 ;
        RECT 88.630 118.215 89.630 118.475 ;
        RECT 89.800 117.820 90.090 118.605 ;
        RECT 90.370 117.820 90.660 138.230 ;
        RECT 87.600 117.530 90.660 117.820 ;
        RECT 91.855 138.230 94.415 138.520 ;
        RECT 91.855 117.820 92.145 138.230 ;
        RECT 92.425 137.435 92.715 138.230 ;
        RECT 92.885 137.575 93.385 137.835 ;
        RECT 92.405 135.405 92.715 137.435 ;
        RECT 92.885 136.295 93.385 136.555 ;
        RECT 93.575 135.405 93.865 138.230 ;
        RECT 92.885 135.015 93.385 135.275 ;
        RECT 92.365 133.015 92.695 134.840 ;
        RECT 93.575 133.015 93.905 134.975 ;
        RECT 92.365 132.725 93.905 133.015 ;
        RECT 92.365 130.890 92.695 132.725 ;
        RECT 93.575 130.890 93.905 132.725 ;
        RECT 92.885 130.455 93.385 130.715 ;
        RECT 92.405 129.445 92.715 130.315 ;
        RECT 93.575 129.445 93.865 130.315 ;
        RECT 92.405 129.165 93.865 129.445 ;
        RECT 92.405 128.285 92.715 129.165 ;
        RECT 92.425 128.165 92.715 128.285 ;
        RECT 93.575 128.165 93.865 129.165 ;
        RECT 92.425 127.885 93.865 128.165 ;
        RECT 92.425 127.755 92.715 127.885 ;
        RECT 92.405 126.885 92.715 127.755 ;
        RECT 93.575 126.885 93.865 127.885 ;
        RECT 92.405 126.605 93.865 126.885 ;
        RECT 92.405 125.725 92.715 126.605 ;
        RECT 93.575 125.725 93.865 126.605 ;
        RECT 92.885 125.335 93.385 125.595 ;
        RECT 93.575 123.490 93.910 125.160 ;
        RECT 92.885 123.055 93.385 123.315 ;
        RECT 93.580 122.880 93.910 123.490 ;
        RECT 93.575 121.210 93.910 122.880 ;
        RECT 92.885 120.775 93.385 121.035 ;
        RECT 92.405 118.605 92.715 120.635 ;
        RECT 92.885 119.495 93.385 119.755 ;
        RECT 92.425 117.820 92.715 118.605 ;
        RECT 92.885 118.215 93.385 118.475 ;
        RECT 93.575 117.820 93.865 120.635 ;
        RECT 94.125 117.820 94.415 138.230 ;
        RECT 91.855 117.530 94.415 117.820 ;
        RECT 80.960 112.980 86.260 113.270 ;
        RECT 88.485 113.280 91.180 113.570 ;
        RECT 91.445 113.280 95.165 113.570 ;
        RECT 63.625 89.140 67.345 89.430 ;
        RECT 67.610 89.140 70.305 89.430 ;
        RECT 88.485 89.430 88.775 113.280 ;
        RECT 89.175 112.625 89.675 112.885 ;
        RECT 89.175 110.345 89.675 110.605 ;
        RECT 89.865 108.500 90.155 113.280 ;
        RECT 92.995 108.500 93.285 113.280 ;
        RECT 93.475 112.625 94.475 112.885 ;
        RECT 93.475 110.345 94.475 110.605 ;
        RECT 89.175 108.065 89.675 108.325 ;
        RECT 93.475 108.065 94.475 108.325 ;
        RECT 89.175 105.785 89.675 106.045 ;
        RECT 89.865 103.940 90.195 107.890 ;
        RECT 90.805 105.775 91.765 106.055 ;
        RECT 89.175 103.505 89.675 103.765 ;
        RECT 91.120 103.330 91.450 105.775 ;
        RECT 92.955 103.940 93.285 107.890 ;
        RECT 93.475 105.785 94.475 106.045 ;
        RECT 93.475 103.505 94.475 103.765 ;
        RECT 89.865 103.000 93.285 103.330 ;
        RECT 89.175 101.225 89.675 101.485 ;
        RECT 89.865 99.380 90.195 103.000 ;
        RECT 90.805 101.215 91.765 101.495 ;
        RECT 89.175 98.945 89.675 99.205 ;
        RECT 91.120 98.770 91.450 101.215 ;
        RECT 92.955 99.380 93.285 103.000 ;
        RECT 93.475 101.225 94.475 101.485 ;
        RECT 93.475 98.945 94.475 99.205 ;
        RECT 89.865 98.440 93.285 98.770 ;
        RECT 89.175 96.665 89.675 96.925 ;
        RECT 89.865 94.820 90.195 98.440 ;
        RECT 92.955 94.820 93.285 98.440 ;
        RECT 93.475 96.665 94.475 96.925 ;
        RECT 89.175 94.385 89.675 94.645 ;
        RECT 93.475 94.385 94.475 94.645 ;
        RECT 89.175 92.105 89.675 92.365 ;
        RECT 89.175 89.825 89.675 90.085 ;
        RECT 89.865 89.430 90.155 94.210 ;
        RECT 92.995 89.430 93.285 94.210 ;
        RECT 93.475 92.105 94.475 92.365 ;
        RECT 93.475 89.825 94.475 90.085 ;
        RECT 94.875 89.430 95.165 113.280 ;
        RECT 96.020 112.230 96.310 151.440 ;
        RECT 97.050 150.785 98.050 151.045 ;
        RECT 97.050 150.005 98.050 150.265 ;
        RECT 98.240 149.660 98.530 151.440 ;
        RECT 97.050 149.225 98.050 149.485 ;
        RECT 96.530 145.100 96.860 149.050 ;
        RECT 97.050 146.945 98.050 147.205 ;
        RECT 97.050 144.665 98.050 144.925 ;
        RECT 98.240 144.160 98.530 144.490 ;
        RECT 97.050 143.870 98.530 144.160 ;
        RECT 98.240 143.380 98.530 143.870 ;
        RECT 97.050 143.090 98.530 143.380 ;
        RECT 98.240 142.600 98.530 143.090 ;
        RECT 97.050 142.310 98.530 142.600 ;
        RECT 98.240 141.980 98.530 142.310 ;
        RECT 97.050 141.545 98.050 141.805 ;
        RECT 96.530 128.300 96.860 141.370 ;
        RECT 98.240 139.700 98.530 141.370 ;
        RECT 97.050 139.265 98.050 139.525 ;
        RECT 98.240 137.420 98.530 139.090 ;
        RECT 97.050 136.985 98.050 137.245 ;
        RECT 98.240 135.140 98.530 136.810 ;
        RECT 97.050 134.705 98.050 134.965 ;
        RECT 98.240 132.860 98.530 134.530 ;
        RECT 97.050 132.425 98.050 132.685 ;
        RECT 98.240 130.580 98.530 132.250 ;
        RECT 100.160 130.580 100.450 151.440 ;
        RECT 100.640 141.545 101.640 141.805 ;
        RECT 100.640 139.265 101.640 139.525 ;
        RECT 100.640 136.985 101.640 137.245 ;
        RECT 100.640 134.705 101.640 134.965 ;
        RECT 100.640 132.425 101.640 132.685 ;
        RECT 97.050 130.145 98.050 130.405 ;
        RECT 100.640 130.145 101.640 130.405 ;
        RECT 98.240 128.300 98.530 129.970 ;
        RECT 97.050 127.865 98.050 128.125 ;
        RECT 100.640 127.865 101.640 128.125 ;
        RECT 96.530 114.620 96.860 127.690 ;
        RECT 98.240 126.020 98.530 127.690 ;
        RECT 101.830 126.020 102.160 129.970 ;
        RECT 97.050 125.585 98.050 125.845 ;
        RECT 100.640 125.585 101.640 125.845 ;
        RECT 98.240 123.740 98.530 125.410 ;
        RECT 97.050 123.305 98.050 123.565 ;
        RECT 98.240 121.460 98.530 123.130 ;
        RECT 97.050 121.025 98.050 121.285 ;
        RECT 98.240 119.180 98.530 120.850 ;
        RECT 97.050 118.745 98.050 119.005 ;
        RECT 98.240 116.900 98.530 118.570 ;
        RECT 97.050 116.465 98.050 116.725 ;
        RECT 98.240 114.620 98.530 116.290 ;
        RECT 97.050 114.185 98.050 114.445 ;
        RECT 97.050 113.405 98.050 113.665 ;
        RECT 97.050 112.625 98.050 112.885 ;
        RECT 98.240 112.230 98.530 114.010 ;
        RECT 100.160 112.230 100.450 125.410 ;
        RECT 100.640 123.305 101.640 123.565 ;
        RECT 100.640 121.025 101.640 121.285 ;
        RECT 100.640 118.745 101.640 119.005 ;
        RECT 100.640 116.465 101.640 116.725 ;
        RECT 100.640 114.185 101.640 114.445 ;
        RECT 102.380 112.230 102.670 151.440 ;
        RECT 96.020 111.940 102.670 112.230 ;
        RECT 88.485 89.140 91.180 89.430 ;
        RECT 91.445 89.140 95.165 89.430 ;
        RECT 88.445 82.960 91.140 83.250 ;
        RECT 91.430 82.960 95.150 83.250 ;
        RECT 71.415 82.610 74.390 82.900 ;
        RECT 74.800 82.610 83.760 82.900 ;
        RECT 84.170 82.610 87.145 82.900 ;
        RECT 71.415 78.120 71.705 82.610 ;
        RECT 72.595 82.200 73.445 82.215 ;
        RECT 72.445 81.970 73.445 82.200 ;
        RECT 72.595 81.955 73.445 81.970 ;
        RECT 71.965 81.360 72.255 81.950 ;
        RECT 72.595 81.770 73.445 81.785 ;
        RECT 72.445 81.540 73.445 81.770 ;
        RECT 72.595 81.525 73.445 81.540 ;
        RECT 73.635 81.360 73.925 82.610 ;
        RECT 72.595 81.340 73.445 81.355 ;
        RECT 72.445 81.110 73.445 81.340 ;
        RECT 72.595 81.095 73.445 81.110 ;
        RECT 71.925 80.500 72.255 81.090 ;
        RECT 72.445 80.665 73.445 80.925 ;
        RECT 73.635 80.500 73.925 81.090 ;
        RECT 72.595 80.480 73.445 80.495 ;
        RECT 72.445 80.250 73.445 80.480 ;
        RECT 72.595 80.235 73.445 80.250 ;
        RECT 71.965 79.640 72.255 80.230 ;
        RECT 73.635 80.100 73.925 80.230 ;
        RECT 74.430 80.100 74.760 82.145 ;
        RECT 75.265 81.360 75.555 82.610 ;
        RECT 75.820 82.200 76.670 82.215 ;
        RECT 77.395 82.200 78.245 82.215 ;
        RECT 75.745 81.970 76.745 82.200 ;
        RECT 77.395 81.970 78.395 82.200 ;
        RECT 75.820 81.955 76.670 81.970 ;
        RECT 77.395 81.955 78.245 81.970 ;
        RECT 78.625 81.950 78.915 82.610 ;
        RECT 75.820 81.770 76.670 81.785 ;
        RECT 77.395 81.770 78.245 81.785 ;
        RECT 75.745 81.540 76.745 81.770 ;
        RECT 77.395 81.540 78.395 81.770 ;
        RECT 75.820 81.525 76.670 81.540 ;
        RECT 77.395 81.525 78.245 81.540 ;
        RECT 78.585 81.360 78.915 81.950 ;
        RECT 75.745 81.095 76.745 81.355 ;
        RECT 77.395 81.340 78.245 81.355 ;
        RECT 77.395 81.110 78.395 81.340 ;
        RECT 77.395 81.095 78.245 81.110 ;
        RECT 75.225 80.100 75.555 81.090 ;
        RECT 75.745 80.665 76.745 80.925 ;
        RECT 77.395 80.665 78.395 80.925 ;
        RECT 75.745 80.235 76.745 80.495 ;
        RECT 77.395 80.480 78.245 80.495 ;
        RECT 77.395 80.250 78.395 80.480 ;
        RECT 77.395 80.235 78.245 80.250 ;
        RECT 72.445 79.805 73.445 80.065 ;
        RECT 73.635 79.770 75.555 80.100 ;
        RECT 75.745 79.805 76.745 80.065 ;
        RECT 77.395 79.805 78.395 80.065 ;
        RECT 73.635 79.640 73.925 79.770 ;
        RECT 75.225 79.640 75.555 79.770 ;
        RECT 78.585 79.640 78.915 81.090 ;
        RECT 72.595 79.620 73.445 79.635 ;
        RECT 72.445 79.390 73.445 79.620 ;
        RECT 72.595 79.375 73.445 79.390 ;
        RECT 75.745 79.375 76.745 79.635 ;
        RECT 77.395 79.620 78.245 79.635 ;
        RECT 77.395 79.390 78.395 79.620 ;
        RECT 77.395 79.375 78.245 79.390 ;
        RECT 71.965 78.780 72.255 79.370 ;
        RECT 72.595 79.190 73.445 79.205 ;
        RECT 72.445 78.960 73.445 79.190 ;
        RECT 72.595 78.945 73.445 78.960 ;
        RECT 72.595 78.760 73.445 78.775 ;
        RECT 72.445 78.530 73.445 78.760 ;
        RECT 72.595 78.515 73.445 78.530 ;
        RECT 72.595 78.120 73.445 78.125 ;
        RECT 73.635 78.120 73.925 79.370 ;
        RECT 75.265 78.120 75.555 79.370 ;
        RECT 75.820 79.190 76.670 79.205 ;
        RECT 77.395 79.190 78.245 79.205 ;
        RECT 75.745 78.960 76.745 79.190 ;
        RECT 77.395 78.960 78.395 79.190 ;
        RECT 75.820 78.945 76.670 78.960 ;
        RECT 77.395 78.945 78.245 78.960 ;
        RECT 78.585 78.780 78.915 79.370 ;
        RECT 75.820 78.760 76.670 78.775 ;
        RECT 77.395 78.760 78.245 78.775 ;
        RECT 75.745 78.530 76.745 78.760 ;
        RECT 77.395 78.530 78.395 78.760 ;
        RECT 75.820 78.515 76.670 78.530 ;
        RECT 77.395 78.515 78.245 78.530 ;
        RECT 75.820 78.120 76.670 78.125 ;
        RECT 77.395 78.120 78.245 78.125 ;
        RECT 78.625 78.120 78.915 78.780 ;
        RECT 79.135 78.120 79.425 82.610 ;
        RECT 79.645 81.950 79.935 82.610 ;
        RECT 80.315 82.200 81.165 82.215 ;
        RECT 81.890 82.200 82.740 82.215 ;
        RECT 80.165 81.970 81.165 82.200 ;
        RECT 81.815 81.970 82.815 82.200 ;
        RECT 80.315 81.955 81.165 81.970 ;
        RECT 81.890 81.955 82.740 81.970 ;
        RECT 79.645 81.360 79.975 81.950 ;
        RECT 80.315 81.770 81.165 81.785 ;
        RECT 81.890 81.770 82.740 81.785 ;
        RECT 80.165 81.540 81.165 81.770 ;
        RECT 81.815 81.540 82.815 81.770 ;
        RECT 80.315 81.525 81.165 81.540 ;
        RECT 81.890 81.525 82.740 81.540 ;
        RECT 83.005 81.360 83.295 82.610 ;
        RECT 80.315 81.340 81.165 81.355 ;
        RECT 80.165 81.110 81.165 81.340 ;
        RECT 80.315 81.095 81.165 81.110 ;
        RECT 81.815 81.095 82.815 81.355 ;
        RECT 79.645 79.640 79.975 81.090 ;
        RECT 80.165 80.665 81.165 80.925 ;
        RECT 81.815 80.665 82.815 80.925 ;
        RECT 80.315 80.480 81.165 80.495 ;
        RECT 80.165 80.250 81.165 80.480 ;
        RECT 80.315 80.235 81.165 80.250 ;
        RECT 81.815 80.235 82.815 80.495 ;
        RECT 83.005 80.100 83.335 81.090 ;
        RECT 83.800 80.100 84.130 82.145 ;
        RECT 84.635 81.360 84.925 82.610 ;
        RECT 85.115 82.200 85.965 82.215 ;
        RECT 85.115 81.970 86.115 82.200 ;
        RECT 85.115 81.955 85.965 81.970 ;
        RECT 85.115 81.770 85.965 81.785 ;
        RECT 85.115 81.540 86.115 81.770 ;
        RECT 85.115 81.525 85.965 81.540 ;
        RECT 86.305 81.360 86.595 81.950 ;
        RECT 85.115 81.340 85.965 81.355 ;
        RECT 85.115 81.110 86.115 81.340 ;
        RECT 85.115 81.095 85.965 81.110 ;
        RECT 84.635 80.500 84.925 81.090 ;
        RECT 85.115 80.665 86.115 80.925 ;
        RECT 86.305 80.500 86.635 81.090 ;
        RECT 85.115 80.480 85.965 80.495 ;
        RECT 85.115 80.250 86.115 80.480 ;
        RECT 85.115 80.235 85.965 80.250 ;
        RECT 84.635 80.100 84.925 80.230 ;
        RECT 80.165 79.805 81.165 80.065 ;
        RECT 81.815 79.805 82.815 80.065 ;
        RECT 83.005 79.770 84.925 80.100 ;
        RECT 85.115 79.805 86.115 80.065 ;
        RECT 83.005 79.640 83.335 79.770 ;
        RECT 84.635 79.640 84.925 79.770 ;
        RECT 86.305 79.640 86.595 80.230 ;
        RECT 80.315 79.620 81.165 79.635 ;
        RECT 80.165 79.390 81.165 79.620 ;
        RECT 80.315 79.375 81.165 79.390 ;
        RECT 81.815 79.375 82.815 79.635 ;
        RECT 85.115 79.620 85.965 79.635 ;
        RECT 85.115 79.390 86.115 79.620 ;
        RECT 85.115 79.375 85.965 79.390 ;
        RECT 79.645 78.780 79.975 79.370 ;
        RECT 80.315 79.190 81.165 79.205 ;
        RECT 81.890 79.190 82.740 79.205 ;
        RECT 80.165 78.960 81.165 79.190 ;
        RECT 81.815 78.960 82.815 79.190 ;
        RECT 80.315 78.945 81.165 78.960 ;
        RECT 81.890 78.945 82.740 78.960 ;
        RECT 79.645 78.120 79.935 78.780 ;
        RECT 80.315 78.760 81.165 78.775 ;
        RECT 81.890 78.760 82.740 78.775 ;
        RECT 80.165 78.530 81.165 78.760 ;
        RECT 81.815 78.530 82.815 78.760 ;
        RECT 80.315 78.515 81.165 78.530 ;
        RECT 81.890 78.515 82.740 78.530 ;
        RECT 80.315 78.120 81.165 78.125 ;
        RECT 81.890 78.120 82.740 78.125 ;
        RECT 83.005 78.120 83.295 79.370 ;
        RECT 84.635 78.120 84.925 79.370 ;
        RECT 85.115 79.190 85.965 79.205 ;
        RECT 85.115 78.960 86.115 79.190 ;
        RECT 85.115 78.945 85.965 78.960 ;
        RECT 86.305 78.780 86.595 79.370 ;
        RECT 85.115 78.760 85.965 78.775 ;
        RECT 85.115 78.530 86.115 78.760 ;
        RECT 85.115 78.515 85.965 78.530 ;
        RECT 85.115 78.120 85.965 78.125 ;
        RECT 86.855 78.120 87.145 82.610 ;
        RECT 88.445 78.470 88.735 82.960 ;
        RECT 89.110 82.305 90.110 82.565 ;
        RECT 89.110 81.875 90.110 82.135 ;
        RECT 90.300 81.710 90.590 82.960 ;
        RECT 89.110 81.445 90.110 81.705 ;
        RECT 89.110 81.015 90.110 81.275 ;
        RECT 90.300 80.880 90.590 81.440 ;
        RECT 91.120 80.880 91.450 82.555 ;
        RECT 91.980 81.710 92.270 82.960 ;
        RECT 92.960 82.550 93.960 82.565 ;
        RECT 92.460 82.320 94.460 82.550 ;
        RECT 92.960 82.305 93.960 82.320 ;
        RECT 92.960 82.120 93.960 82.135 ;
        RECT 92.460 81.890 94.460 82.120 ;
        RECT 92.960 81.875 93.960 81.890 ;
        RECT 92.960 81.690 93.960 81.705 ;
        RECT 92.460 81.460 94.460 81.690 ;
        RECT 92.960 81.445 93.960 81.460 ;
        RECT 91.980 80.880 92.270 81.440 ;
        RECT 92.460 81.015 94.460 81.275 ;
        RECT 89.110 80.585 90.110 80.845 ;
        RECT 90.300 80.550 92.270 80.880 ;
        RECT 92.960 80.830 93.960 80.845 ;
        RECT 92.460 80.600 94.460 80.830 ;
        RECT 92.960 80.585 93.960 80.600 ;
        RECT 89.110 80.155 90.110 80.415 ;
        RECT 90.300 79.990 90.590 80.550 ;
        RECT 91.980 79.990 92.270 80.550 ;
        RECT 92.460 80.155 94.460 80.415 ;
        RECT 89.110 79.725 90.110 79.985 ;
        RECT 92.960 79.970 93.960 79.985 ;
        RECT 92.460 79.740 94.460 79.970 ;
        RECT 92.960 79.725 93.960 79.740 ;
        RECT 89.110 79.295 90.110 79.555 ;
        RECT 89.110 78.865 90.110 79.125 ;
        RECT 90.300 78.470 90.590 79.720 ;
        RECT 91.980 78.470 92.270 79.720 ;
        RECT 92.960 79.540 93.960 79.555 ;
        RECT 92.460 79.310 94.460 79.540 ;
        RECT 92.960 79.295 93.960 79.310 ;
        RECT 92.960 79.110 93.960 79.125 ;
        RECT 92.460 78.880 94.460 79.110 ;
        RECT 92.960 78.865 93.960 78.880 ;
        RECT 94.860 78.470 95.150 82.960 ;
        RECT 88.445 78.180 91.140 78.470 ;
        RECT 91.430 78.180 95.150 78.470 ;
        RECT 71.415 77.830 74.390 78.120 ;
        RECT 74.800 77.830 83.760 78.120 ;
        RECT 84.170 77.830 87.145 78.120 ;
        RECT 64.665 72.300 67.360 72.590 ;
        RECT 67.650 72.300 71.370 72.590 ;
        RECT 64.665 63.510 64.955 72.300 ;
        RECT 65.330 71.645 66.330 71.905 ;
        RECT 65.330 71.215 66.330 71.475 ;
        RECT 66.520 71.050 66.810 72.300 ;
        RECT 65.330 70.785 66.330 71.045 ;
        RECT 65.330 70.355 66.330 70.615 ;
        RECT 66.520 70.235 66.810 70.780 ;
        RECT 67.340 70.235 67.670 71.895 ;
        RECT 68.200 71.050 68.490 72.300 ;
        RECT 69.180 71.890 70.180 71.905 ;
        RECT 68.680 71.660 70.680 71.890 ;
        RECT 69.180 71.645 70.180 71.660 ;
        RECT 69.180 71.460 70.180 71.475 ;
        RECT 68.680 71.230 70.680 71.460 ;
        RECT 69.180 71.215 70.180 71.230 ;
        RECT 69.180 71.030 70.180 71.045 ;
        RECT 68.680 70.800 70.680 71.030 ;
        RECT 69.180 70.785 70.180 70.800 ;
        RECT 68.200 70.235 68.490 70.780 ;
        RECT 68.680 70.355 70.680 70.615 ;
        RECT 65.330 69.925 66.330 70.185 ;
        RECT 66.520 69.905 68.490 70.235 ;
        RECT 69.180 70.170 70.180 70.185 ;
        RECT 68.680 69.940 70.680 70.170 ;
        RECT 69.180 69.925 70.180 69.940 ;
        RECT 65.330 69.495 66.330 69.755 ;
        RECT 66.520 69.330 66.810 69.905 ;
        RECT 67.025 69.485 67.985 69.765 ;
        RECT 65.330 69.065 66.330 69.325 ;
        RECT 65.330 68.635 66.330 68.895 ;
        RECT 65.330 68.205 66.330 68.465 ;
        RECT 65.330 67.775 66.330 68.035 ;
        RECT 65.330 67.345 66.330 67.605 ;
        RECT 66.520 67.210 66.810 69.060 ;
        RECT 67.340 67.210 67.670 69.485 ;
        RECT 68.200 69.330 68.490 69.905 ;
        RECT 68.680 69.495 70.680 69.755 ;
        RECT 69.180 69.310 70.180 69.325 ;
        RECT 68.680 69.080 70.680 69.310 ;
        RECT 69.180 69.065 70.180 69.080 ;
        RECT 68.200 67.210 68.490 69.060 ;
        RECT 68.680 68.635 70.680 68.895 ;
        RECT 69.180 68.450 70.180 68.465 ;
        RECT 68.680 68.220 70.680 68.450 ;
        RECT 69.180 68.205 70.180 68.220 ;
        RECT 68.680 67.775 70.680 68.035 ;
        RECT 69.180 67.590 70.180 67.605 ;
        RECT 68.680 67.360 70.680 67.590 ;
        RECT 69.180 67.345 70.180 67.360 ;
        RECT 65.330 66.915 66.330 67.175 ;
        RECT 66.520 66.880 68.490 67.210 ;
        RECT 68.680 66.915 70.680 67.175 ;
        RECT 65.330 66.485 66.330 66.745 ;
        RECT 65.330 66.055 66.330 66.315 ;
        RECT 65.330 65.625 66.330 65.885 ;
        RECT 65.330 65.195 66.330 65.455 ;
        RECT 66.520 65.030 66.810 66.880 ;
        RECT 68.200 65.030 68.490 66.880 ;
        RECT 69.180 66.730 70.180 66.745 ;
        RECT 68.680 66.500 70.680 66.730 ;
        RECT 69.180 66.485 70.180 66.500 ;
        RECT 68.680 66.055 70.680 66.315 ;
        RECT 69.180 65.870 70.180 65.885 ;
        RECT 68.680 65.640 70.680 65.870 ;
        RECT 69.180 65.625 70.180 65.640 ;
        RECT 68.680 65.195 70.680 65.455 ;
        RECT 65.330 64.765 66.330 65.025 ;
        RECT 69.180 65.010 70.180 65.025 ;
        RECT 68.680 64.780 70.680 65.010 ;
        RECT 69.180 64.765 70.180 64.780 ;
        RECT 65.330 64.335 66.330 64.595 ;
        RECT 65.330 63.905 66.330 64.165 ;
        RECT 66.520 63.510 66.810 64.760 ;
        RECT 68.200 63.510 68.490 64.760 ;
        RECT 69.180 64.580 70.180 64.595 ;
        RECT 68.680 64.350 70.680 64.580 ;
        RECT 69.180 64.335 70.180 64.350 ;
        RECT 69.180 64.150 70.180 64.165 ;
        RECT 68.680 63.920 70.680 64.150 ;
        RECT 69.180 63.905 70.180 63.920 ;
        RECT 71.080 63.510 71.370 72.300 ;
        RECT 64.665 63.220 67.360 63.510 ;
        RECT 67.650 63.220 71.370 63.510 ;
        RECT 73.685 72.300 76.380 72.590 ;
        RECT 76.670 72.300 83.820 72.590 ;
        RECT 84.110 72.300 86.805 72.590 ;
        RECT 73.685 63.510 73.975 72.300 ;
        RECT 74.350 71.645 75.350 71.905 ;
        RECT 74.350 71.215 75.350 71.475 ;
        RECT 75.540 71.050 75.830 72.300 ;
        RECT 74.350 70.785 75.350 71.045 ;
        RECT 74.350 70.355 75.350 70.615 ;
        RECT 75.540 70.235 75.830 70.780 ;
        RECT 76.360 70.235 76.690 71.895 ;
        RECT 77.220 71.050 77.510 72.300 ;
        RECT 78.200 71.890 79.200 71.905 ;
        RECT 77.700 71.660 79.700 71.890 ;
        RECT 78.200 71.645 79.200 71.660 ;
        RECT 78.200 71.460 79.200 71.475 ;
        RECT 77.700 71.230 79.700 71.460 ;
        RECT 78.200 71.215 79.200 71.230 ;
        RECT 78.200 71.030 79.200 71.045 ;
        RECT 77.700 70.800 79.700 71.030 ;
        RECT 78.200 70.785 79.200 70.800 ;
        RECT 77.220 70.235 77.510 70.780 ;
        RECT 77.700 70.355 79.700 70.615 ;
        RECT 74.350 69.925 75.350 70.185 ;
        RECT 75.540 69.905 77.510 70.235 ;
        RECT 78.200 70.170 79.200 70.185 ;
        RECT 77.700 69.940 79.700 70.170 ;
        RECT 78.200 69.925 79.200 69.940 ;
        RECT 74.350 69.495 75.350 69.755 ;
        RECT 75.540 69.330 75.830 69.905 ;
        RECT 76.045 69.485 77.005 69.765 ;
        RECT 74.350 69.065 75.350 69.325 ;
        RECT 74.350 68.635 75.350 68.895 ;
        RECT 74.350 68.205 75.350 68.465 ;
        RECT 74.350 67.775 75.350 68.035 ;
        RECT 74.350 67.345 75.350 67.605 ;
        RECT 75.540 67.210 75.830 69.060 ;
        RECT 76.360 67.210 76.690 69.485 ;
        RECT 77.220 69.330 77.510 69.905 ;
        RECT 77.700 69.495 79.700 69.755 ;
        RECT 78.200 69.310 79.200 69.325 ;
        RECT 77.700 69.080 79.700 69.310 ;
        RECT 78.200 69.065 79.200 69.080 ;
        RECT 77.220 67.210 77.510 69.060 ;
        RECT 77.700 68.635 79.700 68.895 ;
        RECT 78.200 68.450 79.200 68.465 ;
        RECT 77.700 68.220 79.700 68.450 ;
        RECT 78.200 68.205 79.200 68.220 ;
        RECT 77.700 67.775 79.700 68.035 ;
        RECT 78.200 67.590 79.200 67.605 ;
        RECT 77.700 67.360 79.700 67.590 ;
        RECT 78.200 67.345 79.200 67.360 ;
        RECT 74.350 66.915 75.350 67.175 ;
        RECT 75.540 66.880 77.510 67.210 ;
        RECT 77.700 66.915 79.700 67.175 ;
        RECT 74.350 66.485 75.350 66.745 ;
        RECT 74.350 66.055 75.350 66.315 ;
        RECT 74.350 65.625 75.350 65.885 ;
        RECT 74.350 65.195 75.350 65.455 ;
        RECT 75.540 65.030 75.830 66.880 ;
        RECT 77.220 65.030 77.510 66.880 ;
        RECT 78.200 66.730 79.200 66.745 ;
        RECT 77.700 66.500 79.700 66.730 ;
        RECT 78.200 66.485 79.200 66.500 ;
        RECT 77.700 66.055 79.700 66.315 ;
        RECT 78.200 65.870 79.200 65.885 ;
        RECT 77.700 65.640 79.700 65.870 ;
        RECT 78.200 65.625 79.200 65.640 ;
        RECT 77.700 65.195 79.700 65.455 ;
        RECT 74.350 64.765 75.350 65.025 ;
        RECT 78.200 65.010 79.200 65.025 ;
        RECT 77.700 64.780 79.700 65.010 ;
        RECT 78.200 64.765 79.200 64.780 ;
        RECT 74.350 64.335 75.350 64.595 ;
        RECT 74.350 63.905 75.350 64.165 ;
        RECT 75.540 63.510 75.830 64.760 ;
        RECT 77.220 63.510 77.510 64.760 ;
        RECT 78.200 64.580 79.200 64.595 ;
        RECT 77.700 64.350 79.700 64.580 ;
        RECT 78.200 64.335 79.200 64.350 ;
        RECT 78.200 64.150 79.200 64.165 ;
        RECT 77.700 63.920 79.700 64.150 ;
        RECT 78.200 63.905 79.200 63.920 ;
        RECT 80.100 63.510 80.390 72.300 ;
        RECT 81.290 71.890 82.290 71.905 ;
        RECT 80.790 71.660 82.790 71.890 ;
        RECT 81.290 71.645 82.290 71.660 ;
        RECT 81.290 71.460 82.290 71.475 ;
        RECT 80.790 71.230 82.790 71.460 ;
        RECT 81.290 71.215 82.290 71.230 ;
        RECT 82.980 71.050 83.270 72.300 ;
        RECT 81.290 71.030 82.290 71.045 ;
        RECT 80.790 70.800 82.790 71.030 ;
        RECT 81.290 70.785 82.290 70.800 ;
        RECT 80.790 70.355 82.790 70.615 ;
        RECT 82.980 70.235 83.270 70.780 ;
        RECT 83.800 70.235 84.130 71.895 ;
        RECT 84.660 71.050 84.950 72.300 ;
        RECT 85.140 71.645 86.140 71.905 ;
        RECT 85.140 71.215 86.140 71.475 ;
        RECT 85.140 70.785 86.140 71.045 ;
        RECT 84.660 70.235 84.950 70.780 ;
        RECT 85.140 70.355 86.140 70.615 ;
        RECT 81.290 70.170 82.290 70.185 ;
        RECT 80.790 69.940 82.790 70.170 ;
        RECT 81.290 69.925 82.290 69.940 ;
        RECT 82.980 69.905 84.950 70.235 ;
        RECT 85.140 69.925 86.140 70.185 ;
        RECT 80.790 69.495 82.790 69.755 ;
        RECT 82.980 69.330 83.270 69.905 ;
        RECT 83.485 69.485 84.445 69.765 ;
        RECT 81.290 69.310 82.290 69.325 ;
        RECT 80.790 69.080 82.790 69.310 ;
        RECT 81.290 69.065 82.290 69.080 ;
        RECT 80.790 68.635 82.790 68.895 ;
        RECT 81.290 68.450 82.290 68.465 ;
        RECT 80.790 68.220 82.790 68.450 ;
        RECT 81.290 68.205 82.290 68.220 ;
        RECT 80.790 67.775 82.790 68.035 ;
        RECT 81.290 67.590 82.290 67.605 ;
        RECT 80.790 67.360 82.790 67.590 ;
        RECT 81.290 67.345 82.290 67.360 ;
        RECT 82.980 67.210 83.270 69.060 ;
        RECT 83.800 67.210 84.130 69.485 ;
        RECT 84.660 69.330 84.950 69.905 ;
        RECT 85.140 69.495 86.140 69.755 ;
        RECT 85.140 69.065 86.140 69.325 ;
        RECT 84.660 67.210 84.950 69.060 ;
        RECT 85.140 68.635 86.140 68.895 ;
        RECT 85.140 68.205 86.140 68.465 ;
        RECT 85.140 67.775 86.140 68.035 ;
        RECT 85.140 67.345 86.140 67.605 ;
        RECT 80.790 66.915 82.790 67.175 ;
        RECT 82.980 66.880 84.950 67.210 ;
        RECT 85.140 66.915 86.140 67.175 ;
        RECT 81.290 66.730 82.290 66.745 ;
        RECT 80.790 66.500 82.790 66.730 ;
        RECT 81.290 66.485 82.290 66.500 ;
        RECT 80.790 66.055 82.790 66.315 ;
        RECT 81.290 65.870 82.290 65.885 ;
        RECT 80.790 65.640 82.790 65.870 ;
        RECT 81.290 65.625 82.290 65.640 ;
        RECT 80.790 65.195 82.790 65.455 ;
        RECT 82.980 65.030 83.270 66.880 ;
        RECT 84.660 65.030 84.950 66.880 ;
        RECT 85.140 66.485 86.140 66.745 ;
        RECT 85.140 66.055 86.140 66.315 ;
        RECT 85.140 65.625 86.140 65.885 ;
        RECT 85.140 65.195 86.140 65.455 ;
        RECT 81.290 65.010 82.290 65.025 ;
        RECT 80.790 64.780 82.790 65.010 ;
        RECT 81.290 64.765 82.290 64.780 ;
        RECT 85.140 64.765 86.140 65.025 ;
        RECT 81.290 64.580 82.290 64.595 ;
        RECT 80.790 64.350 82.790 64.580 ;
        RECT 81.290 64.335 82.290 64.350 ;
        RECT 81.290 64.150 82.290 64.165 ;
        RECT 80.790 63.920 82.790 64.150 ;
        RECT 81.290 63.905 82.290 63.920 ;
        RECT 82.980 63.510 83.270 64.760 ;
        RECT 84.660 63.510 84.950 64.760 ;
        RECT 85.140 64.335 86.140 64.595 ;
        RECT 85.140 63.905 86.140 64.165 ;
        RECT 86.515 63.510 86.805 72.300 ;
        RECT 73.685 63.220 76.380 63.510 ;
        RECT 76.670 63.220 83.820 63.510 ;
        RECT 84.110 63.220 86.805 63.510 ;
        RECT 88.445 72.300 91.140 72.590 ;
        RECT 91.430 72.300 95.150 72.590 ;
        RECT 88.445 63.510 88.735 72.300 ;
        RECT 89.110 71.645 90.110 71.905 ;
        RECT 89.110 71.215 90.110 71.475 ;
        RECT 90.300 71.050 90.590 72.300 ;
        RECT 89.110 70.785 90.110 71.045 ;
        RECT 89.110 70.355 90.110 70.615 ;
        RECT 90.300 70.235 90.590 70.780 ;
        RECT 91.120 70.235 91.450 71.895 ;
        RECT 91.980 71.050 92.270 72.300 ;
        RECT 92.960 71.890 93.960 71.905 ;
        RECT 92.460 71.660 94.460 71.890 ;
        RECT 92.960 71.645 93.960 71.660 ;
        RECT 92.960 71.460 93.960 71.475 ;
        RECT 92.460 71.230 94.460 71.460 ;
        RECT 92.960 71.215 93.960 71.230 ;
        RECT 92.960 71.030 93.960 71.045 ;
        RECT 92.460 70.800 94.460 71.030 ;
        RECT 92.960 70.785 93.960 70.800 ;
        RECT 91.980 70.235 92.270 70.780 ;
        RECT 92.460 70.355 94.460 70.615 ;
        RECT 89.110 69.925 90.110 70.185 ;
        RECT 90.300 69.905 92.270 70.235 ;
        RECT 92.960 70.170 93.960 70.185 ;
        RECT 92.460 69.940 94.460 70.170 ;
        RECT 92.960 69.925 93.960 69.940 ;
        RECT 89.110 69.495 90.110 69.755 ;
        RECT 90.300 69.330 90.590 69.905 ;
        RECT 90.805 69.485 91.765 69.765 ;
        RECT 89.110 69.065 90.110 69.325 ;
        RECT 89.110 68.635 90.110 68.895 ;
        RECT 89.110 68.205 90.110 68.465 ;
        RECT 89.110 67.775 90.110 68.035 ;
        RECT 89.110 67.345 90.110 67.605 ;
        RECT 90.300 67.210 90.590 69.060 ;
        RECT 91.120 67.210 91.450 69.485 ;
        RECT 91.980 69.330 92.270 69.905 ;
        RECT 92.460 69.495 94.460 69.755 ;
        RECT 92.960 69.310 93.960 69.325 ;
        RECT 92.460 69.080 94.460 69.310 ;
        RECT 92.960 69.065 93.960 69.080 ;
        RECT 91.980 67.210 92.270 69.060 ;
        RECT 92.460 68.635 94.460 68.895 ;
        RECT 92.960 68.450 93.960 68.465 ;
        RECT 92.460 68.220 94.460 68.450 ;
        RECT 92.960 68.205 93.960 68.220 ;
        RECT 92.460 67.775 94.460 68.035 ;
        RECT 92.960 67.590 93.960 67.605 ;
        RECT 92.460 67.360 94.460 67.590 ;
        RECT 92.960 67.345 93.960 67.360 ;
        RECT 89.110 66.915 90.110 67.175 ;
        RECT 90.300 66.880 92.270 67.210 ;
        RECT 92.460 66.915 94.460 67.175 ;
        RECT 89.110 66.485 90.110 66.745 ;
        RECT 89.110 66.055 90.110 66.315 ;
        RECT 89.110 65.625 90.110 65.885 ;
        RECT 89.110 65.195 90.110 65.455 ;
        RECT 90.300 65.030 90.590 66.880 ;
        RECT 91.980 65.030 92.270 66.880 ;
        RECT 92.960 66.730 93.960 66.745 ;
        RECT 92.460 66.500 94.460 66.730 ;
        RECT 92.960 66.485 93.960 66.500 ;
        RECT 92.460 66.055 94.460 66.315 ;
        RECT 92.960 65.870 93.960 65.885 ;
        RECT 92.460 65.640 94.460 65.870 ;
        RECT 92.960 65.625 93.960 65.640 ;
        RECT 92.460 65.195 94.460 65.455 ;
        RECT 89.110 64.765 90.110 65.025 ;
        RECT 92.960 65.010 93.960 65.025 ;
        RECT 92.460 64.780 94.460 65.010 ;
        RECT 92.960 64.765 93.960 64.780 ;
        RECT 89.110 64.335 90.110 64.595 ;
        RECT 89.110 63.905 90.110 64.165 ;
        RECT 90.300 63.510 90.590 64.760 ;
        RECT 91.980 63.510 92.270 64.760 ;
        RECT 92.960 64.580 93.960 64.595 ;
        RECT 92.460 64.350 94.460 64.580 ;
        RECT 92.960 64.335 93.960 64.350 ;
        RECT 92.960 64.150 93.960 64.165 ;
        RECT 92.460 63.920 94.460 64.150 ;
        RECT 92.960 63.905 93.960 63.920 ;
        RECT 94.860 63.510 95.150 72.300 ;
        RECT 88.445 63.220 91.140 63.510 ;
        RECT 91.430 63.220 95.150 63.510 ;
        RECT 108.575 63.320 108.865 164.690 ;
        RECT 109.605 164.035 110.305 164.295 ;
        RECT 109.605 161.755 110.305 162.015 ;
        RECT 110.495 159.910 110.785 164.690 ;
        RECT 110.975 164.035 111.675 164.295 ;
        RECT 110.975 161.755 111.675 162.015 ;
        RECT 111.865 159.910 112.155 164.690 ;
        RECT 112.345 164.035 113.045 164.295 ;
        RECT 112.345 161.755 113.045 162.015 ;
        RECT 109.605 159.475 110.305 159.735 ;
        RECT 110.975 159.475 111.675 159.735 ;
        RECT 112.345 159.475 113.045 159.735 ;
        RECT 110.475 157.465 110.805 159.300 ;
        RECT 111.845 157.465 112.175 159.300 ;
        RECT 109.605 157.185 113.045 157.465 ;
        RECT 109.605 154.915 110.305 155.175 ;
        RECT 110.475 152.905 110.805 157.185 ;
        RECT 110.975 154.915 111.675 155.175 ;
        RECT 111.845 152.905 112.175 157.185 ;
        RECT 112.345 154.915 113.045 155.175 ;
        RECT 109.605 152.625 113.045 152.905 ;
        RECT 109.605 150.355 110.305 150.615 ;
        RECT 110.475 148.345 110.805 152.625 ;
        RECT 110.975 150.355 111.675 150.615 ;
        RECT 111.845 148.345 112.175 152.625 ;
        RECT 112.345 150.355 113.045 150.615 ;
        RECT 109.605 148.065 113.045 148.345 ;
        RECT 109.605 145.795 110.305 146.055 ;
        RECT 110.475 143.785 110.805 148.065 ;
        RECT 110.975 145.795 111.675 146.055 ;
        RECT 111.845 143.785 112.175 148.065 ;
        RECT 112.345 145.795 113.045 146.055 ;
        RECT 109.605 143.505 113.045 143.785 ;
        RECT 109.605 141.235 110.305 141.495 ;
        RECT 110.475 139.225 110.805 143.505 ;
        RECT 110.975 141.235 111.675 141.495 ;
        RECT 111.845 139.225 112.175 143.505 ;
        RECT 112.345 141.235 113.045 141.495 ;
        RECT 109.605 138.945 113.045 139.225 ;
        RECT 109.605 136.675 110.305 136.935 ;
        RECT 109.605 134.395 110.305 134.655 ;
        RECT 109.605 132.115 110.305 132.375 ;
        RECT 109.605 129.835 110.305 130.095 ;
        RECT 109.605 127.555 110.305 127.815 ;
        RECT 109.605 125.275 110.305 125.535 ;
        RECT 109.605 122.995 110.305 123.255 ;
        RECT 109.605 120.715 110.305 120.975 ;
        RECT 109.605 118.435 110.305 118.695 ;
        RECT 109.605 116.155 110.305 116.415 ;
        RECT 109.605 113.875 110.305 114.135 ;
        RECT 109.605 111.595 110.305 111.855 ;
        RECT 109.605 109.315 110.305 109.575 ;
        RECT 109.605 107.035 110.305 107.295 ;
        RECT 109.605 104.755 110.305 105.015 ;
        RECT 109.605 102.475 110.305 102.735 ;
        RECT 109.605 100.195 110.305 100.455 ;
        RECT 109.605 97.915 110.305 98.175 ;
        RECT 109.605 95.635 110.305 95.895 ;
        RECT 109.605 93.355 110.305 93.615 ;
        RECT 109.605 91.075 110.305 91.335 ;
        RECT 109.605 88.795 110.305 89.055 ;
        RECT 109.605 86.515 110.305 86.775 ;
        RECT 109.605 84.235 110.305 84.495 ;
        RECT 109.605 81.955 110.305 82.215 ;
        RECT 109.605 79.675 110.305 79.935 ;
        RECT 109.605 77.395 110.305 77.655 ;
        RECT 109.605 75.115 110.305 75.375 ;
        RECT 109.605 72.835 110.305 73.095 ;
        RECT 109.605 70.555 110.305 70.815 ;
        RECT 110.475 68.710 110.805 138.945 ;
        RECT 110.975 136.675 111.675 136.935 ;
        RECT 110.975 134.395 111.675 134.655 ;
        RECT 110.975 132.115 111.675 132.375 ;
        RECT 110.975 129.835 111.675 130.095 ;
        RECT 110.975 127.555 111.675 127.815 ;
        RECT 110.975 125.275 111.675 125.535 ;
        RECT 110.975 122.995 111.675 123.255 ;
        RECT 110.975 120.715 111.675 120.975 ;
        RECT 110.975 118.435 111.675 118.695 ;
        RECT 110.975 116.155 111.675 116.415 ;
        RECT 110.975 113.875 111.675 114.135 ;
        RECT 110.975 111.595 111.675 111.855 ;
        RECT 110.975 109.315 111.675 109.575 ;
        RECT 110.975 107.035 111.675 107.295 ;
        RECT 110.975 104.755 111.675 105.015 ;
        RECT 110.975 102.475 111.675 102.735 ;
        RECT 110.975 100.195 111.675 100.455 ;
        RECT 110.975 97.915 111.675 98.175 ;
        RECT 110.975 95.635 111.675 95.895 ;
        RECT 110.975 93.355 111.675 93.615 ;
        RECT 110.975 91.075 111.675 91.335 ;
        RECT 110.975 88.795 111.675 89.055 ;
        RECT 110.975 86.515 111.675 86.775 ;
        RECT 110.975 84.235 111.675 84.495 ;
        RECT 110.975 81.955 111.675 82.215 ;
        RECT 110.975 79.675 111.675 79.935 ;
        RECT 110.975 77.395 111.675 77.655 ;
        RECT 110.975 75.115 111.675 75.375 ;
        RECT 110.975 72.835 111.675 73.095 ;
        RECT 110.975 70.555 111.675 70.815 ;
        RECT 111.845 68.710 112.175 138.945 ;
        RECT 112.345 136.675 113.045 136.935 ;
        RECT 112.345 134.395 113.045 134.655 ;
        RECT 112.345 132.115 113.045 132.375 ;
        RECT 112.345 129.835 113.045 130.095 ;
        RECT 112.345 127.555 113.045 127.815 ;
        RECT 112.345 125.275 113.045 125.535 ;
        RECT 112.345 122.995 113.045 123.255 ;
        RECT 112.345 120.715 113.045 120.975 ;
        RECT 112.345 118.435 113.045 118.695 ;
        RECT 112.345 116.155 113.045 116.415 ;
        RECT 112.345 113.875 113.045 114.135 ;
        RECT 113.785 113.755 114.075 164.690 ;
        RECT 121.780 164.650 125.910 164.940 ;
        RECT 114.865 118.095 117.625 118.385 ;
        RECT 114.865 114.545 115.155 118.095 ;
        RECT 116.100 117.725 116.390 118.095 ;
        RECT 115.895 117.495 116.595 117.725 ;
        RECT 115.375 116.180 115.705 117.420 ;
        RECT 116.100 117.295 116.390 117.495 ;
        RECT 115.895 117.065 116.595 117.295 ;
        RECT 116.785 117.065 117.075 118.095 ;
        RECT 115.895 116.620 116.595 116.880 ;
        RECT 115.895 116.190 116.595 116.450 ;
        RECT 115.895 115.760 116.595 116.020 ;
        RECT 115.895 115.345 116.595 115.575 ;
        RECT 116.100 115.145 116.390 115.345 ;
        RECT 115.895 114.915 116.595 115.145 ;
        RECT 116.100 114.545 116.390 114.915 ;
        RECT 116.785 114.545 117.075 115.575 ;
        RECT 117.335 115.090 117.625 118.095 ;
        RECT 118.135 117.860 121.195 118.150 ;
        RECT 118.135 115.090 118.425 117.860 ;
        RECT 118.685 115.110 118.975 117.860 ;
        RECT 119.485 117.490 119.775 117.860 ;
        RECT 119.165 117.260 120.165 117.490 ;
        RECT 119.485 117.060 119.775 117.260 ;
        RECT 119.165 116.830 120.165 117.060 ;
        RECT 119.485 116.630 119.775 116.830 ;
        RECT 119.165 116.400 120.165 116.630 ;
        RECT 119.485 116.200 119.775 116.400 ;
        RECT 119.165 115.970 120.165 116.200 ;
        RECT 119.485 115.770 119.775 115.970 ;
        RECT 119.165 115.540 120.165 115.770 ;
        RECT 119.485 115.340 119.775 115.540 ;
        RECT 120.905 115.435 121.195 117.860 ;
        RECT 121.780 115.435 122.070 164.650 ;
        RECT 122.330 159.910 122.620 164.650 ;
        RECT 122.810 164.035 123.510 164.295 ;
        RECT 122.810 161.755 123.510 162.015 ;
        RECT 122.810 159.475 123.510 159.735 ;
        RECT 122.330 157.630 122.620 159.300 ;
        RECT 122.810 157.195 123.510 157.455 ;
        RECT 122.330 155.350 122.620 157.020 ;
        RECT 122.810 154.915 123.510 155.175 ;
        RECT 122.330 153.070 122.620 154.740 ;
        RECT 122.810 152.635 123.510 152.895 ;
        RECT 122.330 150.790 122.620 152.460 ;
        RECT 122.810 150.355 123.510 150.615 ;
        RECT 122.330 148.510 122.620 150.180 ;
        RECT 122.810 148.075 123.510 148.335 ;
        RECT 122.330 146.230 122.620 147.900 ;
        RECT 122.810 145.795 123.510 146.055 ;
        RECT 122.330 143.950 122.620 145.620 ;
        RECT 122.810 143.515 123.510 143.775 ;
        RECT 122.330 141.670 122.620 143.340 ;
        RECT 122.810 141.235 123.510 141.495 ;
        RECT 122.330 139.390 122.620 141.060 ;
        RECT 122.810 138.955 123.510 139.215 ;
        RECT 122.330 137.110 122.620 138.780 ;
        RECT 122.810 136.675 123.510 136.935 ;
        RECT 122.330 134.830 122.620 136.500 ;
        RECT 122.810 134.395 123.510 134.655 ;
        RECT 122.330 132.550 122.620 134.220 ;
        RECT 122.810 132.115 123.510 132.375 ;
        RECT 122.330 130.270 122.620 131.940 ;
        RECT 122.810 129.835 123.510 130.095 ;
        RECT 122.330 127.990 122.620 129.660 ;
        RECT 122.810 127.555 123.510 127.815 ;
        RECT 122.330 125.710 122.620 127.380 ;
        RECT 122.810 125.275 123.510 125.535 ;
        RECT 122.330 123.430 122.620 125.100 ;
        RECT 122.810 122.995 123.510 123.255 ;
        RECT 122.330 121.150 122.620 122.820 ;
        RECT 122.810 120.715 123.510 120.975 ;
        RECT 122.330 118.870 122.620 120.540 ;
        RECT 122.810 118.435 123.510 118.695 ;
        RECT 122.330 116.590 122.620 118.260 ;
        RECT 122.810 116.155 123.510 116.415 ;
        RECT 119.165 115.110 120.165 115.340 ;
        RECT 117.335 114.545 118.425 115.090 ;
        RECT 119.485 114.910 119.775 115.110 ;
        RECT 119.165 114.680 120.165 114.910 ;
        RECT 114.865 114.255 118.425 114.545 ;
        RECT 118.135 114.050 118.425 114.255 ;
        RECT 119.165 114.235 120.165 114.495 ;
        RECT 118.135 113.820 120.165 114.050 ;
        RECT 113.785 113.465 117.625 113.755 ;
        RECT 112.345 111.595 113.045 111.855 ;
        RECT 113.785 111.635 115.155 113.465 ;
        RECT 115.415 112.395 115.705 113.465 ;
        RECT 116.100 113.055 116.390 113.465 ;
        RECT 115.895 112.825 116.595 113.055 ;
        RECT 116.100 112.625 116.390 112.825 ;
        RECT 115.895 112.395 116.595 112.625 ;
        RECT 115.895 111.950 116.595 112.210 ;
        RECT 112.345 109.315 113.045 109.575 ;
        RECT 112.345 107.035 113.045 107.295 ;
        RECT 112.345 104.755 113.045 105.015 ;
        RECT 112.345 102.475 113.045 102.735 ;
        RECT 112.345 100.195 113.045 100.455 ;
        RECT 112.345 97.915 113.045 98.175 ;
        RECT 112.345 95.635 113.045 95.895 ;
        RECT 112.345 93.355 113.045 93.615 ;
        RECT 112.345 91.075 113.045 91.335 ;
        RECT 112.345 88.795 113.045 89.055 ;
        RECT 112.345 86.515 113.045 86.775 ;
        RECT 112.345 84.235 113.045 84.495 ;
        RECT 112.345 81.955 113.045 82.215 ;
        RECT 112.345 79.675 113.045 79.935 ;
        RECT 113.785 79.555 114.075 111.635 ;
        RECT 114.865 109.835 115.155 111.635 ;
        RECT 115.895 111.520 116.595 111.780 ;
        RECT 115.895 111.090 116.595 111.350 ;
        RECT 115.415 109.835 115.705 110.905 ;
        RECT 115.895 110.675 116.595 110.905 ;
        RECT 116.100 110.475 116.390 110.675 ;
        RECT 115.895 110.245 116.595 110.475 ;
        RECT 116.100 109.835 116.390 110.245 ;
        RECT 116.785 110.120 117.115 111.765 ;
        RECT 117.335 109.835 117.625 113.465 ;
        RECT 114.865 109.545 117.625 109.835 ;
        RECT 118.135 110.010 118.425 113.820 ;
        RECT 119.165 113.375 120.165 113.635 ;
        RECT 120.355 113.390 120.685 114.485 ;
        RECT 120.905 113.435 122.070 115.435 ;
        RECT 122.330 114.310 122.620 115.980 ;
        RECT 122.810 113.875 123.510 114.135 ;
        RECT 119.165 112.960 120.165 113.190 ;
        RECT 119.485 112.760 119.775 112.960 ;
        RECT 118.685 110.010 118.975 112.760 ;
        RECT 119.165 112.530 120.165 112.760 ;
        RECT 119.485 112.330 119.775 112.530 ;
        RECT 119.165 112.100 120.165 112.330 ;
        RECT 119.485 111.900 119.775 112.100 ;
        RECT 119.165 111.670 120.165 111.900 ;
        RECT 119.485 111.470 119.775 111.670 ;
        RECT 119.165 111.240 120.165 111.470 ;
        RECT 119.485 111.040 119.775 111.240 ;
        RECT 119.165 110.810 120.165 111.040 ;
        RECT 119.485 110.610 119.775 110.810 ;
        RECT 119.165 110.380 120.165 110.610 ;
        RECT 119.485 110.010 119.775 110.380 ;
        RECT 120.905 110.010 121.195 113.435 ;
        RECT 118.135 109.720 121.195 110.010 ;
        RECT 114.865 83.895 117.625 84.185 ;
        RECT 114.865 80.345 115.155 83.895 ;
        RECT 116.100 83.525 116.390 83.895 ;
        RECT 115.895 83.295 116.595 83.525 ;
        RECT 115.375 81.980 115.705 83.220 ;
        RECT 116.100 83.095 116.390 83.295 ;
        RECT 115.895 82.865 116.595 83.095 ;
        RECT 116.785 82.865 117.075 83.895 ;
        RECT 115.895 82.420 116.595 82.680 ;
        RECT 115.895 81.990 116.595 82.250 ;
        RECT 115.895 81.560 116.595 81.820 ;
        RECT 115.895 81.145 116.595 81.375 ;
        RECT 116.100 80.945 116.390 81.145 ;
        RECT 115.895 80.715 116.595 80.945 ;
        RECT 116.100 80.345 116.390 80.715 ;
        RECT 116.785 80.345 117.075 81.375 ;
        RECT 117.335 80.890 117.625 83.895 ;
        RECT 118.135 83.660 121.195 83.950 ;
        RECT 118.135 80.890 118.425 83.660 ;
        RECT 118.685 80.910 118.975 83.660 ;
        RECT 119.485 83.290 119.775 83.660 ;
        RECT 119.165 83.060 120.165 83.290 ;
        RECT 119.485 82.860 119.775 83.060 ;
        RECT 119.165 82.630 120.165 82.860 ;
        RECT 119.485 82.430 119.775 82.630 ;
        RECT 119.165 82.200 120.165 82.430 ;
        RECT 119.485 82.000 119.775 82.200 ;
        RECT 119.165 81.770 120.165 82.000 ;
        RECT 119.485 81.570 119.775 81.770 ;
        RECT 119.165 81.340 120.165 81.570 ;
        RECT 119.485 81.140 119.775 81.340 ;
        RECT 119.165 80.910 120.165 81.140 ;
        RECT 117.335 80.345 118.425 80.890 ;
        RECT 119.485 80.710 119.775 80.910 ;
        RECT 119.165 80.480 120.165 80.710 ;
        RECT 114.865 80.055 118.425 80.345 ;
        RECT 118.135 79.850 118.425 80.055 ;
        RECT 119.165 80.035 120.165 80.295 ;
        RECT 118.135 79.620 120.165 79.850 ;
        RECT 113.785 79.265 117.625 79.555 ;
        RECT 112.345 77.395 113.045 77.655 ;
        RECT 113.785 77.435 115.155 79.265 ;
        RECT 115.415 78.195 115.705 79.265 ;
        RECT 116.100 78.855 116.390 79.265 ;
        RECT 115.895 78.625 116.595 78.855 ;
        RECT 116.100 78.425 116.390 78.625 ;
        RECT 115.895 78.195 116.595 78.425 ;
        RECT 115.895 77.750 116.595 78.010 ;
        RECT 112.345 75.115 113.045 75.375 ;
        RECT 112.345 72.835 113.045 73.095 ;
        RECT 112.345 70.555 113.045 70.815 ;
        RECT 109.605 68.275 110.305 68.535 ;
        RECT 110.975 68.275 111.675 68.535 ;
        RECT 112.345 68.275 113.045 68.535 ;
        RECT 109.605 65.995 110.305 66.255 ;
        RECT 109.605 63.715 110.305 63.975 ;
        RECT 110.495 63.320 110.785 68.100 ;
        RECT 110.975 65.995 111.675 66.255 ;
        RECT 110.975 63.715 111.675 63.975 ;
        RECT 111.865 63.320 112.155 68.100 ;
        RECT 112.345 65.995 113.045 66.255 ;
        RECT 112.345 63.715 113.045 63.975 ;
        RECT 113.785 63.320 114.075 77.435 ;
        RECT 114.865 75.635 115.155 77.435 ;
        RECT 115.895 77.320 116.595 77.580 ;
        RECT 115.895 76.890 116.595 77.150 ;
        RECT 115.415 75.635 115.705 76.705 ;
        RECT 115.895 76.475 116.595 76.705 ;
        RECT 116.100 76.275 116.390 76.475 ;
        RECT 115.895 76.045 116.595 76.275 ;
        RECT 116.100 75.635 116.390 76.045 ;
        RECT 116.785 75.920 117.115 77.565 ;
        RECT 117.335 75.635 117.625 79.265 ;
        RECT 114.865 75.345 117.625 75.635 ;
        RECT 118.135 75.810 118.425 79.620 ;
        RECT 119.165 79.175 120.165 79.435 ;
        RECT 120.355 79.190 120.685 80.285 ;
        RECT 120.905 79.435 121.195 83.660 ;
        RECT 121.780 79.435 122.070 113.435 ;
        RECT 122.330 112.030 122.620 113.700 ;
        RECT 122.810 111.595 123.510 111.855 ;
        RECT 122.330 109.750 122.620 111.420 ;
        RECT 122.810 109.315 123.510 109.575 ;
        RECT 122.330 107.470 122.620 109.140 ;
        RECT 122.810 107.035 123.510 107.295 ;
        RECT 122.330 105.190 122.620 106.860 ;
        RECT 122.810 104.755 123.510 105.015 ;
        RECT 122.330 102.910 122.620 104.580 ;
        RECT 122.810 102.475 123.510 102.735 ;
        RECT 122.330 100.630 122.620 102.300 ;
        RECT 122.810 100.195 123.510 100.455 ;
        RECT 122.330 98.350 122.620 100.020 ;
        RECT 122.810 97.915 123.510 98.175 ;
        RECT 122.330 96.070 122.620 97.740 ;
        RECT 122.810 95.635 123.510 95.895 ;
        RECT 122.330 93.790 122.620 95.460 ;
        RECT 122.810 93.355 123.510 93.615 ;
        RECT 122.330 91.510 122.620 93.180 ;
        RECT 122.810 91.075 123.510 91.335 ;
        RECT 122.330 89.040 122.620 90.900 ;
        RECT 122.810 89.040 123.510 89.055 ;
        RECT 122.330 88.810 123.510 89.040 ;
        RECT 122.330 86.760 122.620 88.810 ;
        RECT 122.810 88.795 123.510 88.810 ;
        RECT 122.810 86.760 123.510 86.775 ;
        RECT 122.330 86.530 123.510 86.760 ;
        RECT 122.330 84.670 122.620 86.530 ;
        RECT 122.810 86.515 123.510 86.530 ;
        RECT 122.810 84.235 123.510 84.495 ;
        RECT 122.330 80.110 122.620 84.060 ;
        RECT 123.680 82.770 124.010 164.160 ;
        RECT 124.180 164.035 124.880 164.295 ;
        RECT 124.180 161.755 124.880 162.015 ;
        RECT 125.070 159.910 125.360 164.650 ;
        RECT 124.180 159.475 124.880 159.735 ;
        RECT 125.070 157.630 125.360 159.300 ;
        RECT 124.180 157.195 124.880 157.455 ;
        RECT 125.070 155.350 125.360 157.020 ;
        RECT 124.180 154.915 124.880 155.175 ;
        RECT 125.070 153.070 125.360 154.740 ;
        RECT 124.180 152.635 124.880 152.895 ;
        RECT 125.070 150.790 125.360 152.460 ;
        RECT 124.180 150.355 124.880 150.615 ;
        RECT 125.070 148.510 125.360 150.180 ;
        RECT 124.180 148.075 124.880 148.335 ;
        RECT 125.070 146.230 125.360 147.900 ;
        RECT 124.180 145.795 124.880 146.055 ;
        RECT 125.070 143.950 125.360 145.620 ;
        RECT 124.180 143.515 124.880 143.775 ;
        RECT 125.070 141.670 125.360 143.340 ;
        RECT 124.180 141.235 124.880 141.495 ;
        RECT 125.070 139.390 125.360 141.060 ;
        RECT 124.180 138.955 124.880 139.215 ;
        RECT 125.070 137.110 125.360 138.780 ;
        RECT 124.180 136.675 124.880 136.935 ;
        RECT 125.070 134.830 125.360 136.500 ;
        RECT 124.180 134.395 124.880 134.655 ;
        RECT 125.070 132.550 125.360 134.220 ;
        RECT 124.180 132.115 124.880 132.375 ;
        RECT 125.070 130.270 125.360 131.940 ;
        RECT 124.180 129.835 124.880 130.095 ;
        RECT 125.070 127.990 125.360 129.660 ;
        RECT 124.180 127.555 124.880 127.815 ;
        RECT 125.070 125.710 125.360 127.380 ;
        RECT 124.180 125.275 124.880 125.535 ;
        RECT 125.070 123.430 125.360 125.100 ;
        RECT 124.180 122.995 124.880 123.255 ;
        RECT 125.070 121.150 125.360 122.820 ;
        RECT 124.180 120.715 124.880 120.975 ;
        RECT 125.070 118.870 125.360 120.540 ;
        RECT 124.180 118.435 124.880 118.695 ;
        RECT 125.070 116.590 125.360 118.260 ;
        RECT 124.180 116.155 124.880 116.415 ;
        RECT 125.070 114.310 125.360 115.980 ;
        RECT 124.180 113.875 124.880 114.135 ;
        RECT 125.070 112.030 125.360 113.700 ;
        RECT 124.180 111.595 124.880 111.855 ;
        RECT 125.070 109.750 125.360 111.420 ;
        RECT 124.180 109.315 124.880 109.575 ;
        RECT 125.070 107.470 125.360 109.140 ;
        RECT 124.180 107.035 124.880 107.295 ;
        RECT 125.070 105.190 125.360 106.860 ;
        RECT 124.180 104.755 124.880 105.015 ;
        RECT 125.070 102.910 125.360 104.580 ;
        RECT 124.180 102.475 124.880 102.735 ;
        RECT 125.070 100.630 125.360 102.300 ;
        RECT 124.180 100.195 124.880 100.455 ;
        RECT 125.070 98.350 125.360 100.020 ;
        RECT 124.180 97.915 124.880 98.175 ;
        RECT 125.070 96.070 125.360 97.740 ;
        RECT 124.180 95.635 124.880 95.895 ;
        RECT 125.070 93.790 125.360 95.460 ;
        RECT 124.180 93.355 124.880 93.615 ;
        RECT 125.070 91.510 125.360 93.180 ;
        RECT 124.180 91.075 124.880 91.335 ;
        RECT 124.180 89.040 124.880 89.055 ;
        RECT 125.070 89.040 125.360 90.900 ;
        RECT 124.180 88.810 125.360 89.040 ;
        RECT 124.180 88.795 124.880 88.810 ;
        RECT 124.180 86.760 124.880 86.775 ;
        RECT 125.070 86.760 125.360 88.810 ;
        RECT 124.180 86.530 125.360 86.760 ;
        RECT 124.180 86.515 124.880 86.530 ;
        RECT 124.180 84.480 124.880 84.495 ;
        RECT 125.070 84.480 125.360 86.530 ;
        RECT 124.180 84.250 125.360 84.480 ;
        RECT 124.180 84.235 124.880 84.250 ;
        RECT 122.810 81.955 123.510 82.215 ;
        RECT 124.180 82.200 124.880 82.215 ;
        RECT 125.070 82.200 125.360 84.250 ;
        RECT 124.180 81.970 125.360 82.200 ;
        RECT 124.180 81.955 124.880 81.970 ;
        RECT 122.810 79.675 123.510 79.935 ;
        RECT 124.180 79.675 124.880 79.935 ;
        RECT 119.165 78.760 120.165 78.990 ;
        RECT 119.485 78.560 119.775 78.760 ;
        RECT 118.685 75.810 118.975 78.560 ;
        RECT 119.165 78.330 120.165 78.560 ;
        RECT 119.485 78.130 119.775 78.330 ;
        RECT 119.165 77.900 120.165 78.130 ;
        RECT 119.485 77.700 119.775 77.900 ;
        RECT 119.165 77.470 120.165 77.700 ;
        RECT 119.485 77.270 119.775 77.470 ;
        RECT 120.905 77.435 122.070 79.435 ;
        RECT 119.165 77.040 120.165 77.270 ;
        RECT 119.485 76.840 119.775 77.040 ;
        RECT 119.165 76.610 120.165 76.840 ;
        RECT 119.485 76.410 119.775 76.610 ;
        RECT 119.165 76.180 120.165 76.410 ;
        RECT 119.485 75.810 119.775 76.180 ;
        RECT 120.905 75.810 121.195 77.435 ;
        RECT 121.780 77.040 122.070 77.435 ;
        RECT 122.330 77.040 122.620 79.500 ;
        RECT 122.810 77.395 123.510 77.655 ;
        RECT 123.700 77.040 123.990 79.500 ;
        RECT 124.180 77.395 124.880 77.655 ;
        RECT 125.070 77.040 125.360 81.970 ;
        RECT 125.620 77.040 125.910 164.650 ;
        RECT 121.780 76.750 125.910 77.040 ;
        RECT 118.135 75.520 121.195 75.810 ;
        RECT 108.575 63.030 114.075 63.320 ;
        RECT 114.715 70.580 117.475 70.860 ;
        RECT 114.715 70.570 123.885 70.580 ;
        RECT 114.715 60.400 115.005 70.570 ;
        RECT 115.745 69.915 116.445 70.175 ;
        RECT 115.225 63.510 115.555 69.690 ;
        RECT 116.635 68.070 116.925 70.570 ;
        RECT 117.185 70.290 123.885 70.570 ;
        RECT 117.185 68.060 118.700 70.290 ;
        RECT 118.960 69.220 119.250 70.290 ;
        RECT 119.440 69.635 120.140 69.895 ;
        RECT 119.440 69.205 120.140 69.465 ;
        RECT 119.440 68.775 120.140 69.035 ;
        RECT 119.440 68.360 120.140 68.620 ;
        RECT 115.745 67.635 116.445 67.895 ;
        RECT 115.745 65.355 116.445 65.615 ;
        RECT 115.745 63.075 116.445 63.335 ;
        RECT 115.745 60.795 116.445 61.055 ;
        RECT 116.635 60.400 116.925 62.900 ;
        RECT 117.185 60.400 117.475 68.060 ;
        RECT 118.410 65.800 118.700 68.060 ;
        RECT 119.440 67.915 120.140 68.175 ;
        RECT 119.440 67.500 120.140 67.760 ;
        RECT 120.330 67.500 120.660 69.980 ;
        RECT 121.675 69.220 121.965 70.290 ;
        RECT 122.360 69.880 122.650 70.290 ;
        RECT 122.155 69.650 122.855 69.880 ;
        RECT 122.360 69.450 122.650 69.650 ;
        RECT 122.155 69.220 122.855 69.450 ;
        RECT 122.155 68.775 122.855 69.035 ;
        RECT 122.155 68.345 122.855 68.605 ;
        RECT 122.155 67.915 122.855 68.175 ;
        RECT 122.155 67.485 122.855 67.745 ;
        RECT 123.045 67.500 123.375 70.055 ;
        RECT 119.440 67.055 120.140 67.315 ;
        RECT 122.155 67.055 122.855 67.315 ;
        RECT 118.960 65.800 119.250 66.870 ;
        RECT 119.440 66.625 120.140 66.885 ;
        RECT 119.440 66.195 120.140 66.455 ;
        RECT 121.675 65.800 121.965 66.870 ;
        RECT 122.155 66.640 122.855 66.870 ;
        RECT 122.360 66.440 122.650 66.640 ;
        RECT 122.155 66.210 122.855 66.440 ;
        RECT 122.360 65.800 122.650 66.210 ;
        RECT 123.595 65.800 123.885 70.290 ;
        RECT 118.410 65.510 123.885 65.800 ;
        RECT 124.395 70.250 127.155 70.540 ;
        RECT 114.715 60.110 117.475 60.400 ;
        RECT 118.410 65.000 123.885 65.290 ;
        RECT 118.410 60.590 118.700 65.000 ;
        RECT 118.960 63.970 119.250 65.000 ;
        RECT 119.440 64.385 120.140 64.645 ;
        RECT 119.440 63.955 120.140 64.215 ;
        RECT 119.440 63.525 120.140 63.785 ;
        RECT 120.330 63.625 120.770 64.715 ;
        RECT 121.675 63.970 121.965 65.000 ;
        RECT 122.360 64.630 122.650 65.000 ;
        RECT 122.155 64.400 122.855 64.630 ;
        RECT 122.360 64.200 122.650 64.400 ;
        RECT 122.155 63.970 122.855 64.200 ;
        RECT 119.440 63.110 120.140 63.370 ;
        RECT 119.440 62.665 120.140 62.925 ;
        RECT 119.440 62.250 120.140 62.510 ;
        RECT 120.330 62.250 120.660 63.625 ;
        RECT 122.155 63.525 122.855 63.785 ;
        RECT 123.595 63.365 123.885 65.000 ;
        RECT 124.395 63.365 124.685 70.250 ;
        RECT 124.945 66.640 125.235 70.250 ;
        RECT 125.425 69.635 126.125 69.895 ;
        RECT 125.425 69.205 126.125 69.465 ;
        RECT 125.425 68.775 126.125 69.035 ;
        RECT 125.425 68.345 126.125 68.605 ;
        RECT 125.425 67.915 126.125 68.175 ;
        RECT 125.425 67.485 126.125 67.745 ;
        RECT 125.425 67.055 126.125 67.315 ;
        RECT 125.425 66.625 126.125 66.885 ;
        RECT 125.425 66.195 126.125 66.455 ;
        RECT 125.425 65.765 126.125 66.025 ;
        RECT 125.425 65.335 126.125 65.595 ;
        RECT 125.425 64.905 126.125 65.165 ;
        RECT 126.315 64.920 126.610 66.010 ;
        RECT 125.425 64.475 126.125 64.735 ;
        RECT 122.155 63.095 122.855 63.355 ;
        RECT 122.155 62.665 122.855 62.925 ;
        RECT 122.155 62.235 122.855 62.495 ;
        RECT 119.440 61.805 120.140 62.065 ;
        RECT 122.155 61.805 122.855 62.065 ;
        RECT 118.960 60.590 119.250 61.620 ;
        RECT 119.440 61.375 120.140 61.635 ;
        RECT 119.440 60.945 120.140 61.205 ;
        RECT 121.675 60.590 121.965 61.620 ;
        RECT 122.155 61.390 122.855 61.620 ;
        RECT 122.360 61.190 122.650 61.390 ;
        RECT 122.155 60.960 122.855 61.190 ;
        RECT 122.360 60.590 122.650 60.960 ;
        RECT 123.045 60.935 123.375 63.340 ;
        RECT 123.595 62.225 124.685 63.365 ;
        RECT 123.595 60.590 123.885 62.225 ;
        RECT 118.410 60.300 123.885 60.590 ;
        RECT 124.395 60.680 124.685 62.225 ;
        RECT 124.945 60.680 125.235 64.290 ;
        RECT 125.425 64.045 126.125 64.305 ;
        RECT 125.425 63.615 126.125 63.875 ;
        RECT 125.425 63.185 126.125 63.445 ;
        RECT 125.425 62.755 126.125 63.015 ;
        RECT 125.425 62.325 126.125 62.585 ;
        RECT 125.425 61.895 126.125 62.155 ;
        RECT 125.425 61.465 126.125 61.725 ;
        RECT 125.425 61.035 126.125 61.295 ;
        RECT 126.865 60.680 127.155 70.250 ;
        RECT 124.395 60.390 127.155 60.680 ;
      LAYER via ;
        RECT 108.245 173.855 108.505 174.115 ;
        RECT 108.565 173.855 108.825 174.115 ;
        RECT 108.885 173.855 109.145 174.115 ;
        RECT 112.095 173.855 112.355 174.115 ;
        RECT 112.415 173.855 112.675 174.115 ;
        RECT 112.735 173.855 112.995 174.115 ;
        RECT 108.245 173.185 108.505 173.445 ;
        RECT 108.565 173.185 108.825 173.445 ;
        RECT 108.885 173.185 109.145 173.445 ;
        RECT 108.245 172.755 108.505 173.015 ;
        RECT 108.565 172.755 108.825 173.015 ;
        RECT 108.885 172.755 109.145 173.015 ;
        RECT 110.240 173.090 110.500 173.350 ;
        RECT 110.240 172.770 110.500 173.030 ;
        RECT 108.245 172.325 108.505 172.585 ;
        RECT 108.565 172.325 108.825 172.585 ;
        RECT 108.885 172.325 109.145 172.585 ;
        RECT 108.245 171.895 108.505 172.155 ;
        RECT 108.565 171.895 108.825 172.155 ;
        RECT 108.885 171.895 109.145 172.155 ;
        RECT 112.095 173.185 112.355 173.445 ;
        RECT 112.415 173.185 112.675 173.445 ;
        RECT 112.735 173.185 112.995 173.445 ;
        RECT 112.095 172.755 112.355 173.015 ;
        RECT 112.415 172.755 112.675 173.015 ;
        RECT 112.735 172.755 112.995 173.015 ;
        RECT 112.095 172.325 112.355 172.585 ;
        RECT 112.415 172.325 112.675 172.585 ;
        RECT 112.735 172.325 112.995 172.585 ;
        RECT 111.615 171.895 111.875 172.155 ;
        RECT 111.935 171.895 112.195 172.155 ;
        RECT 112.255 171.895 112.515 172.155 ;
        RECT 112.575 171.895 112.835 172.155 ;
        RECT 112.895 171.895 113.155 172.155 ;
        RECT 113.215 171.895 113.475 172.155 ;
        RECT 108.245 171.465 108.505 171.725 ;
        RECT 108.565 171.465 108.825 171.725 ;
        RECT 108.885 171.465 109.145 171.725 ;
        RECT 112.095 171.465 112.355 171.725 ;
        RECT 112.415 171.465 112.675 171.725 ;
        RECT 112.735 171.465 112.995 171.725 ;
        RECT 108.245 171.035 108.505 171.295 ;
        RECT 108.565 171.035 108.825 171.295 ;
        RECT 108.885 171.035 109.145 171.295 ;
        RECT 111.615 171.035 111.875 171.295 ;
        RECT 111.935 171.035 112.195 171.295 ;
        RECT 112.255 171.035 112.515 171.295 ;
        RECT 112.575 171.035 112.835 171.295 ;
        RECT 112.895 171.035 113.155 171.295 ;
        RECT 113.215 171.035 113.475 171.295 ;
        RECT 108.245 170.605 108.505 170.865 ;
        RECT 108.565 170.605 108.825 170.865 ;
        RECT 108.885 170.605 109.145 170.865 ;
        RECT 112.095 170.605 112.355 170.865 ;
        RECT 112.415 170.605 112.675 170.865 ;
        RECT 112.735 170.605 112.995 170.865 ;
        RECT 108.245 170.175 108.505 170.435 ;
        RECT 108.565 170.175 108.825 170.435 ;
        RECT 108.885 170.175 109.145 170.435 ;
        RECT 108.245 169.745 108.505 170.005 ;
        RECT 108.565 169.745 108.825 170.005 ;
        RECT 108.885 169.745 109.145 170.005 ;
        RECT 112.095 170.175 112.355 170.435 ;
        RECT 112.415 170.175 112.675 170.435 ;
        RECT 112.735 170.175 112.995 170.435 ;
        RECT 112.095 169.745 112.355 170.005 ;
        RECT 112.415 169.745 112.675 170.005 ;
        RECT 112.735 169.745 112.995 170.005 ;
        RECT 108.245 169.075 108.505 169.335 ;
        RECT 108.565 169.075 108.825 169.335 ;
        RECT 108.885 169.075 109.145 169.335 ;
        RECT 112.095 169.075 112.355 169.335 ;
        RECT 112.415 169.075 112.675 169.335 ;
        RECT 112.735 169.075 112.995 169.335 ;
        RECT 109.665 164.705 109.925 164.965 ;
        RECT 109.985 164.705 110.245 164.965 ;
        RECT 111.035 164.705 111.295 164.965 ;
        RECT 111.355 164.705 111.615 164.965 ;
        RECT 112.405 164.705 112.665 164.965 ;
        RECT 112.725 164.705 112.985 164.965 ;
        RECT 57.200 151.455 57.460 151.715 ;
        RECT 57.520 151.455 57.780 151.715 ;
        RECT 57.840 151.455 58.100 151.715 ;
        RECT 60.790 151.455 61.050 151.715 ;
        RECT 61.110 151.455 61.370 151.715 ;
        RECT 61.430 151.455 61.690 151.715 ;
        RECT 57.200 141.545 57.460 141.805 ;
        RECT 57.520 141.545 57.780 141.805 ;
        RECT 57.840 141.545 58.100 141.805 ;
        RECT 57.200 139.265 57.460 139.525 ;
        RECT 57.520 139.265 57.780 139.525 ;
        RECT 57.840 139.265 58.100 139.525 ;
        RECT 57.200 136.985 57.460 137.245 ;
        RECT 57.520 136.985 57.780 137.245 ;
        RECT 57.840 136.985 58.100 137.245 ;
        RECT 57.200 134.705 57.460 134.965 ;
        RECT 57.520 134.705 57.780 134.965 ;
        RECT 57.840 134.705 58.100 134.965 ;
        RECT 57.200 132.425 57.460 132.685 ;
        RECT 57.520 132.425 57.780 132.685 ;
        RECT 57.840 132.425 58.100 132.685 ;
        RECT 60.790 150.785 61.050 151.045 ;
        RECT 61.110 150.785 61.370 151.045 ;
        RECT 61.430 150.785 61.690 151.045 ;
        RECT 60.790 150.005 61.050 150.265 ;
        RECT 61.110 150.005 61.370 150.265 ;
        RECT 61.430 150.005 61.690 150.265 ;
        RECT 60.790 149.225 61.050 149.485 ;
        RECT 61.110 149.225 61.370 149.485 ;
        RECT 61.430 149.225 61.690 149.485 ;
        RECT 61.965 148.790 62.225 149.050 ;
        RECT 61.965 148.470 62.225 148.730 ;
        RECT 61.965 148.150 62.225 148.410 ;
        RECT 60.790 146.945 61.050 147.205 ;
        RECT 61.110 146.945 61.370 147.205 ;
        RECT 61.430 146.945 61.690 147.205 ;
        RECT 60.790 144.665 61.050 144.925 ;
        RECT 61.110 144.665 61.370 144.925 ;
        RECT 61.430 144.665 61.690 144.925 ;
        RECT 60.790 143.885 61.050 144.145 ;
        RECT 61.110 143.885 61.370 144.145 ;
        RECT 61.430 143.885 61.690 144.145 ;
        RECT 60.790 143.105 61.050 143.365 ;
        RECT 61.110 143.105 61.370 143.365 ;
        RECT 61.430 143.105 61.690 143.365 ;
        RECT 60.790 142.325 61.050 142.585 ;
        RECT 61.110 142.325 61.370 142.585 ;
        RECT 61.430 142.325 61.690 142.585 ;
        RECT 60.790 141.545 61.050 141.805 ;
        RECT 61.110 141.545 61.370 141.805 ;
        RECT 61.430 141.545 61.690 141.805 ;
        RECT 61.965 141.110 62.225 141.370 ;
        RECT 61.965 140.790 62.225 141.050 ;
        RECT 61.965 140.470 62.225 140.730 ;
        RECT 60.790 139.265 61.050 139.525 ;
        RECT 61.110 139.265 61.370 139.525 ;
        RECT 61.430 139.265 61.690 139.525 ;
        RECT 60.790 136.985 61.050 137.245 ;
        RECT 61.110 136.985 61.370 137.245 ;
        RECT 61.430 136.985 61.690 137.245 ;
        RECT 60.790 134.705 61.050 134.965 ;
        RECT 61.110 134.705 61.370 134.965 ;
        RECT 61.430 134.705 61.690 134.965 ;
        RECT 60.790 132.425 61.050 132.685 ;
        RECT 61.110 132.425 61.370 132.685 ;
        RECT 61.430 132.425 61.690 132.685 ;
        RECT 57.200 130.145 57.460 130.405 ;
        RECT 57.520 130.145 57.780 130.405 ;
        RECT 57.840 130.145 58.100 130.405 ;
        RECT 60.790 130.145 61.050 130.405 ;
        RECT 61.110 130.145 61.370 130.405 ;
        RECT 61.430 130.145 61.690 130.405 ;
        RECT 56.665 128.185 56.925 128.445 ;
        RECT 56.665 127.865 56.925 128.125 ;
        RECT 57.200 127.865 57.460 128.125 ;
        RECT 57.520 127.865 57.780 128.125 ;
        RECT 57.840 127.865 58.100 128.125 ;
        RECT 60.790 127.865 61.050 128.125 ;
        RECT 61.110 127.865 61.370 128.125 ;
        RECT 61.430 127.865 61.690 128.125 ;
        RECT 56.665 127.545 56.925 127.805 ;
        RECT 57.200 125.585 57.460 125.845 ;
        RECT 57.520 125.585 57.780 125.845 ;
        RECT 57.840 125.585 58.100 125.845 ;
        RECT 60.790 125.585 61.050 125.845 ;
        RECT 61.110 125.585 61.370 125.845 ;
        RECT 61.430 125.585 61.690 125.845 ;
        RECT 57.200 123.305 57.460 123.565 ;
        RECT 57.520 123.305 57.780 123.565 ;
        RECT 57.840 123.305 58.100 123.565 ;
        RECT 57.200 121.025 57.460 121.285 ;
        RECT 57.520 121.025 57.780 121.285 ;
        RECT 57.840 121.025 58.100 121.285 ;
        RECT 57.200 118.745 57.460 119.005 ;
        RECT 57.520 118.745 57.780 119.005 ;
        RECT 57.840 118.745 58.100 119.005 ;
        RECT 57.200 116.465 57.460 116.725 ;
        RECT 57.520 116.465 57.780 116.725 ;
        RECT 57.840 116.465 58.100 116.725 ;
        RECT 57.200 114.185 57.460 114.445 ;
        RECT 57.520 114.185 57.780 114.445 ;
        RECT 57.840 114.185 58.100 114.445 ;
        RECT 60.790 123.305 61.050 123.565 ;
        RECT 61.110 123.305 61.370 123.565 ;
        RECT 61.430 123.305 61.690 123.565 ;
        RECT 60.790 121.025 61.050 121.285 ;
        RECT 61.110 121.025 61.370 121.285 ;
        RECT 61.430 121.025 61.690 121.285 ;
        RECT 60.790 118.745 61.050 119.005 ;
        RECT 61.110 118.745 61.370 119.005 ;
        RECT 61.430 118.745 61.690 119.005 ;
        RECT 60.790 116.465 61.050 116.725 ;
        RECT 61.110 116.465 61.370 116.725 ;
        RECT 61.430 116.465 61.690 116.725 ;
        RECT 61.965 115.260 62.225 115.520 ;
        RECT 61.965 114.940 62.225 115.200 ;
        RECT 61.965 114.620 62.225 114.880 ;
        RECT 60.790 114.185 61.050 114.445 ;
        RECT 61.110 114.185 61.370 114.445 ;
        RECT 61.430 114.185 61.690 114.445 ;
        RECT 60.790 113.405 61.050 113.665 ;
        RECT 61.110 113.405 61.370 113.665 ;
        RECT 61.430 113.405 61.690 113.665 ;
        RECT 60.790 112.625 61.050 112.885 ;
        RECT 61.110 112.625 61.370 112.885 ;
        RECT 61.430 112.625 61.690 112.885 ;
        RECT 65.525 151.455 65.785 151.715 ;
        RECT 65.525 150.785 65.785 151.045 ;
        RECT 65.525 150.005 65.785 150.265 ;
        RECT 65.525 149.225 65.785 149.485 ;
        RECT 64.920 147.265 65.180 147.525 ;
        RECT 64.920 146.945 65.180 147.205 ;
        RECT 65.525 146.945 65.785 147.205 ;
        RECT 64.920 146.625 65.180 146.885 ;
        RECT 65.525 144.665 65.785 144.925 ;
        RECT 65.525 143.885 65.785 144.145 ;
        RECT 65.525 143.105 65.785 143.365 ;
        RECT 93.005 151.455 93.265 151.715 ;
        RECT 65.525 142.435 65.785 142.695 ;
        RECT 73.680 142.735 73.940 142.995 ;
        RECT 76.420 142.735 76.680 142.995 ;
        RECT 65.525 138.245 65.785 138.505 ;
        RECT 65.525 137.575 65.785 137.835 ;
        RECT 65.525 136.295 65.785 136.555 ;
        RECT 65.525 135.015 65.785 135.275 ;
        RECT 64.920 134.715 65.180 134.975 ;
        RECT 64.920 134.395 65.180 134.655 ;
        RECT 64.920 134.075 65.180 134.335 ;
        RECT 66.130 134.580 66.390 134.840 ;
        RECT 66.130 134.260 66.390 134.520 ;
        RECT 66.130 133.940 66.390 134.200 ;
        RECT 65.525 130.455 65.785 130.715 ;
        RECT 65.525 129.175 65.785 129.435 ;
        RECT 65.525 127.895 65.785 128.155 ;
        RECT 65.525 126.615 65.785 126.875 ;
        RECT 65.525 125.335 65.785 125.595 ;
        RECT 64.915 123.375 65.175 123.635 ;
        RECT 64.915 123.055 65.175 123.315 ;
        RECT 65.525 123.055 65.785 123.315 ;
        RECT 64.915 122.735 65.175 122.995 ;
        RECT 65.525 120.775 65.785 121.035 ;
        RECT 65.525 119.495 65.785 119.755 ;
        RECT 65.525 118.215 65.785 118.475 ;
        RECT 65.525 117.545 65.785 117.805 ;
        RECT 69.210 138.245 69.470 138.505 ;
        RECT 69.530 138.245 69.790 138.505 ;
        RECT 69.850 138.245 70.110 138.505 ;
        RECT 69.210 137.575 69.470 137.835 ;
        RECT 69.530 137.575 69.790 137.835 ;
        RECT 69.850 137.575 70.110 137.835 ;
        RECT 69.210 136.295 69.470 136.555 ;
        RECT 69.530 136.295 69.790 136.555 ;
        RECT 69.850 136.295 70.110 136.555 ;
        RECT 69.210 135.015 69.470 135.275 ;
        RECT 69.530 135.015 69.790 135.275 ;
        RECT 69.850 135.015 70.110 135.275 ;
        RECT 69.210 132.715 69.470 132.975 ;
        RECT 69.530 132.715 69.790 132.975 ;
        RECT 69.850 132.715 70.110 132.975 ;
        RECT 68.675 131.530 68.935 131.790 ;
        RECT 68.675 131.210 68.935 131.470 ;
        RECT 68.675 130.890 68.935 131.150 ;
        RECT 69.210 130.455 69.470 130.715 ;
        RECT 69.530 130.455 69.790 130.715 ;
        RECT 69.850 130.455 70.110 130.715 ;
        RECT 69.210 129.175 69.470 129.435 ;
        RECT 69.530 129.175 69.790 129.435 ;
        RECT 69.850 129.175 70.110 129.435 ;
        RECT 69.210 127.895 69.470 128.155 ;
        RECT 69.530 127.895 69.790 128.155 ;
        RECT 69.850 127.895 70.110 128.155 ;
        RECT 69.210 126.615 69.470 126.875 ;
        RECT 69.530 126.615 69.790 126.875 ;
        RECT 69.850 126.615 70.110 126.875 ;
        RECT 69.210 125.335 69.470 125.595 ;
        RECT 69.530 125.335 69.790 125.595 ;
        RECT 69.850 125.335 70.110 125.595 ;
        RECT 69.210 123.025 69.470 123.285 ;
        RECT 69.530 123.025 69.790 123.285 ;
        RECT 69.850 123.025 70.110 123.285 ;
        RECT 69.210 120.775 69.470 121.035 ;
        RECT 69.530 120.775 69.790 121.035 ;
        RECT 69.850 120.775 70.110 121.035 ;
        RECT 69.210 119.495 69.470 119.755 ;
        RECT 69.530 119.495 69.790 119.755 ;
        RECT 69.850 119.495 70.110 119.755 ;
        RECT 69.210 118.215 69.470 118.475 ;
        RECT 69.530 118.215 69.790 118.475 ;
        RECT 69.850 118.215 70.110 118.475 ;
        RECT 69.210 117.545 69.470 117.805 ;
        RECT 69.530 117.545 69.790 117.805 ;
        RECT 69.850 117.545 70.110 117.805 ;
        RECT 57.200 111.955 57.460 112.215 ;
        RECT 57.520 111.955 57.780 112.215 ;
        RECT 57.840 111.955 58.100 112.215 ;
        RECT 60.790 111.955 61.050 112.215 ;
        RECT 61.110 111.955 61.370 112.215 ;
        RECT 61.430 111.955 61.690 112.215 ;
        RECT 64.365 113.295 64.625 113.555 ;
        RECT 64.685 113.295 64.945 113.555 ;
        RECT 65.005 113.295 65.265 113.555 ;
        RECT 69.235 113.295 69.495 113.555 ;
        RECT 64.365 112.625 64.625 112.885 ;
        RECT 64.685 112.625 64.945 112.885 ;
        RECT 65.005 112.625 65.265 112.885 ;
        RECT 64.365 110.345 64.625 110.605 ;
        RECT 64.685 110.345 64.945 110.605 ;
        RECT 65.005 110.345 65.265 110.605 ;
        RECT 69.235 112.625 69.495 112.885 ;
        RECT 69.235 110.345 69.495 110.605 ;
        RECT 64.365 108.065 64.625 108.325 ;
        RECT 64.685 108.065 64.945 108.325 ;
        RECT 65.005 108.065 65.265 108.325 ;
        RECT 69.235 108.065 69.495 108.325 ;
        RECT 65.540 107.630 65.800 107.890 ;
        RECT 65.540 107.310 65.800 107.570 ;
        RECT 65.540 106.990 65.800 107.250 ;
        RECT 64.365 105.785 64.625 106.045 ;
        RECT 64.685 105.785 64.945 106.045 ;
        RECT 65.005 105.785 65.265 106.045 ;
        RECT 68.630 107.630 68.890 107.890 ;
        RECT 68.630 107.310 68.890 107.570 ;
        RECT 68.630 106.990 68.890 107.250 ;
        RECT 67.055 105.785 67.315 106.045 ;
        RECT 67.375 105.785 67.635 106.045 ;
        RECT 67.695 105.785 67.955 106.045 ;
        RECT 64.365 103.505 64.625 103.765 ;
        RECT 64.685 103.505 64.945 103.765 ;
        RECT 65.005 103.505 65.265 103.765 ;
        RECT 69.235 105.785 69.495 106.045 ;
        RECT 69.235 103.505 69.495 103.765 ;
        RECT 64.365 101.225 64.625 101.485 ;
        RECT 64.685 101.225 64.945 101.485 ;
        RECT 65.005 101.225 65.265 101.485 ;
        RECT 67.055 101.225 67.315 101.485 ;
        RECT 67.375 101.225 67.635 101.485 ;
        RECT 67.695 101.225 67.955 101.485 ;
        RECT 64.365 98.945 64.625 99.205 ;
        RECT 64.685 98.945 64.945 99.205 ;
        RECT 65.005 98.945 65.265 99.205 ;
        RECT 69.235 101.225 69.495 101.485 ;
        RECT 69.235 98.945 69.495 99.205 ;
        RECT 64.365 96.665 64.625 96.925 ;
        RECT 64.685 96.665 64.945 96.925 ;
        RECT 65.005 96.665 65.265 96.925 ;
        RECT 69.235 96.665 69.495 96.925 ;
        RECT 64.365 94.385 64.625 94.645 ;
        RECT 64.685 94.385 64.945 94.645 ;
        RECT 65.005 94.385 65.265 94.645 ;
        RECT 69.235 94.385 69.495 94.645 ;
        RECT 64.365 92.105 64.625 92.365 ;
        RECT 64.685 92.105 64.945 92.365 ;
        RECT 65.005 92.105 65.265 92.365 ;
        RECT 64.365 89.825 64.625 90.085 ;
        RECT 64.685 89.825 64.945 90.085 ;
        RECT 65.005 89.825 65.265 90.085 ;
        RECT 69.235 92.105 69.495 92.365 ;
        RECT 69.235 89.825 69.495 90.085 ;
        RECT 73.680 142.105 73.940 142.365 ;
        RECT 73.075 141.110 73.335 141.370 ;
        RECT 73.075 140.790 73.335 141.050 ;
        RECT 73.680 139.545 73.940 139.805 ;
        RECT 73.680 137.265 73.940 137.525 ;
        RECT 76.420 141.705 76.680 141.965 ;
        RECT 76.420 138.425 76.680 138.685 ;
        RECT 73.680 134.985 73.940 135.245 ;
        RECT 76.420 135.145 76.680 135.405 ;
        RECT 73.680 132.705 73.940 132.965 ;
        RECT 73.680 130.425 73.940 130.685 ;
        RECT 73.680 129.145 73.940 129.405 ;
        RECT 73.680 127.865 73.940 128.125 ;
        RECT 76.420 127.865 76.680 128.125 ;
        RECT 73.680 126.585 73.940 126.845 ;
        RECT 77.025 126.785 77.285 127.045 ;
        RECT 77.025 126.465 77.285 126.725 ;
        RECT 77.025 126.145 77.285 126.405 ;
        RECT 77.025 125.825 77.285 126.085 ;
        RECT 73.680 125.305 73.940 125.565 ;
        RECT 73.680 123.025 73.940 123.285 ;
        RECT 73.680 120.745 73.940 121.005 ;
        RECT 76.420 120.585 76.680 120.845 ;
        RECT 73.680 118.465 73.940 118.725 ;
        RECT 73.680 116.185 73.940 116.445 ;
        RECT 73.075 114.940 73.335 115.200 ;
        RECT 73.075 114.620 73.335 114.880 ;
        RECT 73.680 113.625 73.940 113.885 ;
        RECT 76.420 117.305 76.680 117.565 ;
        RECT 76.420 114.025 76.680 114.285 ;
        RECT 73.680 112.995 73.940 113.255 ;
        RECT 76.420 112.995 76.680 113.255 ;
        RECT 82.110 142.735 82.370 142.995 ;
        RECT 84.850 142.735 85.110 142.995 ;
        RECT 82.110 141.705 82.370 141.965 ;
        RECT 82.110 138.425 82.370 138.685 ;
        RECT 84.850 142.105 85.110 142.365 ;
        RECT 85.455 141.110 85.715 141.370 ;
        RECT 85.455 140.790 85.715 141.050 ;
        RECT 84.850 139.545 85.110 139.805 ;
        RECT 84.850 137.265 85.110 137.525 ;
        RECT 82.110 135.145 82.370 135.405 ;
        RECT 84.850 134.985 85.110 135.245 ;
        RECT 84.850 132.705 85.110 132.965 ;
        RECT 84.850 130.425 85.110 130.685 ;
        RECT 84.850 129.145 85.110 129.405 ;
        RECT 82.110 127.865 82.370 128.125 ;
        RECT 84.850 127.865 85.110 128.125 ;
        RECT 81.505 126.785 81.765 127.045 ;
        RECT 81.505 126.465 81.765 126.725 ;
        RECT 81.505 126.145 81.765 126.405 ;
        RECT 81.505 125.825 81.765 126.085 ;
        RECT 84.850 126.585 85.110 126.845 ;
        RECT 84.850 125.305 85.110 125.565 ;
        RECT 84.850 123.025 85.110 123.285 ;
        RECT 82.110 120.585 82.370 120.845 ;
        RECT 84.850 120.745 85.110 121.005 ;
        RECT 82.110 117.305 82.370 117.565 ;
        RECT 82.110 114.025 82.370 114.285 ;
        RECT 84.850 118.465 85.110 118.725 ;
        RECT 84.850 116.185 85.110 116.445 ;
        RECT 85.455 114.940 85.715 115.200 ;
        RECT 85.455 114.620 85.715 114.880 ;
        RECT 84.850 113.625 85.110 113.885 ;
        RECT 93.005 150.785 93.265 151.045 ;
        RECT 93.005 150.005 93.265 150.265 ;
        RECT 93.005 149.225 93.265 149.485 ;
        RECT 93.610 147.265 93.870 147.525 ;
        RECT 93.005 146.945 93.265 147.205 ;
        RECT 93.610 146.945 93.870 147.205 ;
        RECT 93.610 146.625 93.870 146.885 ;
        RECT 93.005 144.665 93.265 144.925 ;
        RECT 93.005 143.885 93.265 144.145 ;
        RECT 93.005 143.105 93.265 143.365 ;
        RECT 93.005 142.435 93.265 142.695 ;
        RECT 97.100 151.455 97.360 151.715 ;
        RECT 97.420 151.455 97.680 151.715 ;
        RECT 97.740 151.455 98.000 151.715 ;
        RECT 100.690 151.455 100.950 151.715 ;
        RECT 101.010 151.455 101.270 151.715 ;
        RECT 101.330 151.455 101.590 151.715 ;
        RECT 88.680 138.245 88.940 138.505 ;
        RECT 89.000 138.245 89.260 138.505 ;
        RECT 89.320 138.245 89.580 138.505 ;
        RECT 88.680 137.575 88.940 137.835 ;
        RECT 89.000 137.575 89.260 137.835 ;
        RECT 89.320 137.575 89.580 137.835 ;
        RECT 88.680 136.295 88.940 136.555 ;
        RECT 89.000 136.295 89.260 136.555 ;
        RECT 89.320 136.295 89.580 136.555 ;
        RECT 88.680 135.015 88.940 135.275 ;
        RECT 89.000 135.015 89.260 135.275 ;
        RECT 89.320 135.015 89.580 135.275 ;
        RECT 88.680 132.715 88.940 132.975 ;
        RECT 89.000 132.715 89.260 132.975 ;
        RECT 89.320 132.715 89.580 132.975 ;
        RECT 89.855 131.530 90.115 131.790 ;
        RECT 89.855 131.210 90.115 131.470 ;
        RECT 89.855 130.890 90.115 131.150 ;
        RECT 88.680 130.455 88.940 130.715 ;
        RECT 89.000 130.455 89.260 130.715 ;
        RECT 89.320 130.455 89.580 130.715 ;
        RECT 88.680 129.175 88.940 129.435 ;
        RECT 89.000 129.175 89.260 129.435 ;
        RECT 89.320 129.175 89.580 129.435 ;
        RECT 88.680 127.895 88.940 128.155 ;
        RECT 89.000 127.895 89.260 128.155 ;
        RECT 89.320 127.895 89.580 128.155 ;
        RECT 88.680 126.615 88.940 126.875 ;
        RECT 89.000 126.615 89.260 126.875 ;
        RECT 89.320 126.615 89.580 126.875 ;
        RECT 88.680 125.335 88.940 125.595 ;
        RECT 89.000 125.335 89.260 125.595 ;
        RECT 89.320 125.335 89.580 125.595 ;
        RECT 88.680 123.025 88.940 123.285 ;
        RECT 89.000 123.025 89.260 123.285 ;
        RECT 89.320 123.025 89.580 123.285 ;
        RECT 88.680 120.775 88.940 121.035 ;
        RECT 89.000 120.775 89.260 121.035 ;
        RECT 89.320 120.775 89.580 121.035 ;
        RECT 88.680 119.495 88.940 119.755 ;
        RECT 89.000 119.495 89.260 119.755 ;
        RECT 89.320 119.495 89.580 119.755 ;
        RECT 88.680 118.215 88.940 118.475 ;
        RECT 89.000 118.215 89.260 118.475 ;
        RECT 89.320 118.215 89.580 118.475 ;
        RECT 88.680 117.545 88.940 117.805 ;
        RECT 89.000 117.545 89.260 117.805 ;
        RECT 89.320 117.545 89.580 117.805 ;
        RECT 93.005 138.245 93.265 138.505 ;
        RECT 93.005 137.575 93.265 137.835 ;
        RECT 93.005 136.295 93.265 136.555 ;
        RECT 93.005 135.015 93.265 135.275 ;
        RECT 92.400 134.580 92.660 134.840 ;
        RECT 92.400 134.260 92.660 134.520 ;
        RECT 92.400 133.940 92.660 134.200 ;
        RECT 93.610 134.715 93.870 134.975 ;
        RECT 93.610 134.395 93.870 134.655 ;
        RECT 93.610 134.075 93.870 134.335 ;
        RECT 93.005 130.455 93.265 130.715 ;
        RECT 93.005 129.175 93.265 129.435 ;
        RECT 93.005 127.895 93.265 128.155 ;
        RECT 93.005 126.615 93.265 126.875 ;
        RECT 93.005 125.335 93.265 125.595 ;
        RECT 93.615 123.375 93.875 123.635 ;
        RECT 93.005 123.055 93.265 123.315 ;
        RECT 93.615 123.055 93.875 123.315 ;
        RECT 93.615 122.735 93.875 122.995 ;
        RECT 93.005 120.775 93.265 121.035 ;
        RECT 93.005 119.495 93.265 119.755 ;
        RECT 93.005 118.215 93.265 118.475 ;
        RECT 93.005 117.545 93.265 117.805 ;
        RECT 82.110 112.995 82.370 113.255 ;
        RECT 84.850 112.995 85.110 113.255 ;
        RECT 89.295 113.295 89.555 113.555 ;
        RECT 93.525 113.295 93.785 113.555 ;
        RECT 93.845 113.295 94.105 113.555 ;
        RECT 94.165 113.295 94.425 113.555 ;
        RECT 64.365 89.155 64.625 89.415 ;
        RECT 64.685 89.155 64.945 89.415 ;
        RECT 65.005 89.155 65.265 89.415 ;
        RECT 69.235 89.155 69.495 89.415 ;
        RECT 89.295 112.625 89.555 112.885 ;
        RECT 89.295 110.345 89.555 110.605 ;
        RECT 93.525 112.625 93.785 112.885 ;
        RECT 93.845 112.625 94.105 112.885 ;
        RECT 94.165 112.625 94.425 112.885 ;
        RECT 93.525 110.345 93.785 110.605 ;
        RECT 93.845 110.345 94.105 110.605 ;
        RECT 94.165 110.345 94.425 110.605 ;
        RECT 89.295 108.065 89.555 108.325 ;
        RECT 93.525 108.065 93.785 108.325 ;
        RECT 93.845 108.065 94.105 108.325 ;
        RECT 94.165 108.065 94.425 108.325 ;
        RECT 89.900 107.630 90.160 107.890 ;
        RECT 89.900 107.310 90.160 107.570 ;
        RECT 89.900 106.990 90.160 107.250 ;
        RECT 89.295 105.785 89.555 106.045 ;
        RECT 92.990 107.630 93.250 107.890 ;
        RECT 92.990 107.310 93.250 107.570 ;
        RECT 92.990 106.990 93.250 107.250 ;
        RECT 90.835 105.785 91.095 106.045 ;
        RECT 91.155 105.785 91.415 106.045 ;
        RECT 91.475 105.785 91.735 106.045 ;
        RECT 89.295 103.505 89.555 103.765 ;
        RECT 93.525 105.785 93.785 106.045 ;
        RECT 93.845 105.785 94.105 106.045 ;
        RECT 94.165 105.785 94.425 106.045 ;
        RECT 93.525 103.505 93.785 103.765 ;
        RECT 93.845 103.505 94.105 103.765 ;
        RECT 94.165 103.505 94.425 103.765 ;
        RECT 89.295 101.225 89.555 101.485 ;
        RECT 90.835 101.225 91.095 101.485 ;
        RECT 91.155 101.225 91.415 101.485 ;
        RECT 91.475 101.225 91.735 101.485 ;
        RECT 89.295 98.945 89.555 99.205 ;
        RECT 93.525 101.225 93.785 101.485 ;
        RECT 93.845 101.225 94.105 101.485 ;
        RECT 94.165 101.225 94.425 101.485 ;
        RECT 93.525 98.945 93.785 99.205 ;
        RECT 93.845 98.945 94.105 99.205 ;
        RECT 94.165 98.945 94.425 99.205 ;
        RECT 89.295 96.665 89.555 96.925 ;
        RECT 93.525 96.665 93.785 96.925 ;
        RECT 93.845 96.665 94.105 96.925 ;
        RECT 94.165 96.665 94.425 96.925 ;
        RECT 89.295 94.385 89.555 94.645 ;
        RECT 93.525 94.385 93.785 94.645 ;
        RECT 93.845 94.385 94.105 94.645 ;
        RECT 94.165 94.385 94.425 94.645 ;
        RECT 89.295 92.105 89.555 92.365 ;
        RECT 89.295 89.825 89.555 90.085 ;
        RECT 93.525 92.105 93.785 92.365 ;
        RECT 93.845 92.105 94.105 92.365 ;
        RECT 94.165 92.105 94.425 92.365 ;
        RECT 93.525 89.825 93.785 90.085 ;
        RECT 93.845 89.825 94.105 90.085 ;
        RECT 94.165 89.825 94.425 90.085 ;
        RECT 97.100 150.785 97.360 151.045 ;
        RECT 97.420 150.785 97.680 151.045 ;
        RECT 97.740 150.785 98.000 151.045 ;
        RECT 97.100 150.005 97.360 150.265 ;
        RECT 97.420 150.005 97.680 150.265 ;
        RECT 97.740 150.005 98.000 150.265 ;
        RECT 97.100 149.225 97.360 149.485 ;
        RECT 97.420 149.225 97.680 149.485 ;
        RECT 97.740 149.225 98.000 149.485 ;
        RECT 96.565 148.790 96.825 149.050 ;
        RECT 96.565 148.470 96.825 148.730 ;
        RECT 96.565 148.150 96.825 148.410 ;
        RECT 97.100 146.945 97.360 147.205 ;
        RECT 97.420 146.945 97.680 147.205 ;
        RECT 97.740 146.945 98.000 147.205 ;
        RECT 97.100 144.665 97.360 144.925 ;
        RECT 97.420 144.665 97.680 144.925 ;
        RECT 97.740 144.665 98.000 144.925 ;
        RECT 97.100 143.885 97.360 144.145 ;
        RECT 97.420 143.885 97.680 144.145 ;
        RECT 97.740 143.885 98.000 144.145 ;
        RECT 97.100 143.105 97.360 143.365 ;
        RECT 97.420 143.105 97.680 143.365 ;
        RECT 97.740 143.105 98.000 143.365 ;
        RECT 97.100 142.325 97.360 142.585 ;
        RECT 97.420 142.325 97.680 142.585 ;
        RECT 97.740 142.325 98.000 142.585 ;
        RECT 97.100 141.545 97.360 141.805 ;
        RECT 97.420 141.545 97.680 141.805 ;
        RECT 97.740 141.545 98.000 141.805 ;
        RECT 96.565 141.110 96.825 141.370 ;
        RECT 96.565 140.790 96.825 141.050 ;
        RECT 96.565 140.470 96.825 140.730 ;
        RECT 97.100 139.265 97.360 139.525 ;
        RECT 97.420 139.265 97.680 139.525 ;
        RECT 97.740 139.265 98.000 139.525 ;
        RECT 97.100 136.985 97.360 137.245 ;
        RECT 97.420 136.985 97.680 137.245 ;
        RECT 97.740 136.985 98.000 137.245 ;
        RECT 97.100 134.705 97.360 134.965 ;
        RECT 97.420 134.705 97.680 134.965 ;
        RECT 97.740 134.705 98.000 134.965 ;
        RECT 97.100 132.425 97.360 132.685 ;
        RECT 97.420 132.425 97.680 132.685 ;
        RECT 97.740 132.425 98.000 132.685 ;
        RECT 100.690 141.545 100.950 141.805 ;
        RECT 101.010 141.545 101.270 141.805 ;
        RECT 101.330 141.545 101.590 141.805 ;
        RECT 100.690 139.265 100.950 139.525 ;
        RECT 101.010 139.265 101.270 139.525 ;
        RECT 101.330 139.265 101.590 139.525 ;
        RECT 100.690 136.985 100.950 137.245 ;
        RECT 101.010 136.985 101.270 137.245 ;
        RECT 101.330 136.985 101.590 137.245 ;
        RECT 100.690 134.705 100.950 134.965 ;
        RECT 101.010 134.705 101.270 134.965 ;
        RECT 101.330 134.705 101.590 134.965 ;
        RECT 100.690 132.425 100.950 132.685 ;
        RECT 101.010 132.425 101.270 132.685 ;
        RECT 101.330 132.425 101.590 132.685 ;
        RECT 97.100 130.145 97.360 130.405 ;
        RECT 97.420 130.145 97.680 130.405 ;
        RECT 97.740 130.145 98.000 130.405 ;
        RECT 100.690 130.145 100.950 130.405 ;
        RECT 101.010 130.145 101.270 130.405 ;
        RECT 101.330 130.145 101.590 130.405 ;
        RECT 101.865 128.185 102.125 128.445 ;
        RECT 97.100 127.865 97.360 128.125 ;
        RECT 97.420 127.865 97.680 128.125 ;
        RECT 97.740 127.865 98.000 128.125 ;
        RECT 100.690 127.865 100.950 128.125 ;
        RECT 101.010 127.865 101.270 128.125 ;
        RECT 101.330 127.865 101.590 128.125 ;
        RECT 101.865 127.865 102.125 128.125 ;
        RECT 101.865 127.545 102.125 127.805 ;
        RECT 97.100 125.585 97.360 125.845 ;
        RECT 97.420 125.585 97.680 125.845 ;
        RECT 97.740 125.585 98.000 125.845 ;
        RECT 100.690 125.585 100.950 125.845 ;
        RECT 101.010 125.585 101.270 125.845 ;
        RECT 101.330 125.585 101.590 125.845 ;
        RECT 97.100 123.305 97.360 123.565 ;
        RECT 97.420 123.305 97.680 123.565 ;
        RECT 97.740 123.305 98.000 123.565 ;
        RECT 97.100 121.025 97.360 121.285 ;
        RECT 97.420 121.025 97.680 121.285 ;
        RECT 97.740 121.025 98.000 121.285 ;
        RECT 97.100 118.745 97.360 119.005 ;
        RECT 97.420 118.745 97.680 119.005 ;
        RECT 97.740 118.745 98.000 119.005 ;
        RECT 97.100 116.465 97.360 116.725 ;
        RECT 97.420 116.465 97.680 116.725 ;
        RECT 97.740 116.465 98.000 116.725 ;
        RECT 96.565 115.260 96.825 115.520 ;
        RECT 96.565 114.940 96.825 115.200 ;
        RECT 96.565 114.620 96.825 114.880 ;
        RECT 97.100 114.185 97.360 114.445 ;
        RECT 97.420 114.185 97.680 114.445 ;
        RECT 97.740 114.185 98.000 114.445 ;
        RECT 97.100 113.405 97.360 113.665 ;
        RECT 97.420 113.405 97.680 113.665 ;
        RECT 97.740 113.405 98.000 113.665 ;
        RECT 97.100 112.625 97.360 112.885 ;
        RECT 97.420 112.625 97.680 112.885 ;
        RECT 97.740 112.625 98.000 112.885 ;
        RECT 100.690 123.305 100.950 123.565 ;
        RECT 101.010 123.305 101.270 123.565 ;
        RECT 101.330 123.305 101.590 123.565 ;
        RECT 100.690 121.025 100.950 121.285 ;
        RECT 101.010 121.025 101.270 121.285 ;
        RECT 101.330 121.025 101.590 121.285 ;
        RECT 100.690 118.745 100.950 119.005 ;
        RECT 101.010 118.745 101.270 119.005 ;
        RECT 101.330 118.745 101.590 119.005 ;
        RECT 100.690 116.465 100.950 116.725 ;
        RECT 101.010 116.465 101.270 116.725 ;
        RECT 101.330 116.465 101.590 116.725 ;
        RECT 100.690 114.185 100.950 114.445 ;
        RECT 101.010 114.185 101.270 114.445 ;
        RECT 101.330 114.185 101.590 114.445 ;
        RECT 97.100 111.955 97.360 112.215 ;
        RECT 97.420 111.955 97.680 112.215 ;
        RECT 97.740 111.955 98.000 112.215 ;
        RECT 100.690 111.955 100.950 112.215 ;
        RECT 101.010 111.955 101.270 112.215 ;
        RECT 101.330 111.955 101.590 112.215 ;
        RECT 89.295 89.155 89.555 89.415 ;
        RECT 93.525 89.155 93.785 89.415 ;
        RECT 93.845 89.155 94.105 89.415 ;
        RECT 94.165 89.155 94.425 89.415 ;
        RECT 89.160 82.975 89.420 83.235 ;
        RECT 89.480 82.975 89.740 83.235 ;
        RECT 89.800 82.975 90.060 83.235 ;
        RECT 93.010 82.975 93.270 83.235 ;
        RECT 93.330 82.975 93.590 83.235 ;
        RECT 93.650 82.975 93.910 83.235 ;
        RECT 72.730 82.625 72.990 82.885 ;
        RECT 73.050 82.625 73.310 82.885 ;
        RECT 75.955 82.625 76.215 82.885 ;
        RECT 76.275 82.625 76.535 82.885 ;
        RECT 77.530 82.625 77.790 82.885 ;
        RECT 77.850 82.625 78.110 82.885 ;
        RECT 80.450 82.625 80.710 82.885 ;
        RECT 80.770 82.625 81.030 82.885 ;
        RECT 82.025 82.625 82.285 82.885 ;
        RECT 82.345 82.625 82.605 82.885 ;
        RECT 85.250 82.625 85.510 82.885 ;
        RECT 85.570 82.625 85.830 82.885 ;
        RECT 72.730 81.955 72.990 82.215 ;
        RECT 73.050 81.955 73.310 82.215 ;
        RECT 72.730 81.525 72.990 81.785 ;
        RECT 73.050 81.525 73.310 81.785 ;
        RECT 74.465 81.745 74.725 82.005 ;
        RECT 74.465 81.425 74.725 81.685 ;
        RECT 72.730 81.095 72.990 81.355 ;
        RECT 73.050 81.095 73.310 81.355 ;
        RECT 71.960 80.825 72.220 81.085 ;
        RECT 71.960 80.505 72.220 80.765 ;
        RECT 72.495 80.665 72.755 80.925 ;
        RECT 72.815 80.665 73.075 80.925 ;
        RECT 73.135 80.665 73.395 80.925 ;
        RECT 72.730 80.235 72.990 80.495 ;
        RECT 73.050 80.235 73.310 80.495 ;
        RECT 75.955 81.955 76.215 82.215 ;
        RECT 76.275 81.955 76.535 82.215 ;
        RECT 77.530 81.955 77.790 82.215 ;
        RECT 77.850 81.955 78.110 82.215 ;
        RECT 75.955 81.525 76.215 81.785 ;
        RECT 76.275 81.525 76.535 81.785 ;
        RECT 77.530 81.525 77.790 81.785 ;
        RECT 77.850 81.525 78.110 81.785 ;
        RECT 75.795 81.095 76.055 81.355 ;
        RECT 76.115 81.095 76.375 81.355 ;
        RECT 76.435 81.095 76.695 81.355 ;
        RECT 77.530 81.095 77.790 81.355 ;
        RECT 77.850 81.095 78.110 81.355 ;
        RECT 75.795 80.665 76.055 80.925 ;
        RECT 76.115 80.665 76.375 80.925 ;
        RECT 76.435 80.665 76.695 80.925 ;
        RECT 77.445 80.665 77.705 80.925 ;
        RECT 77.765 80.665 78.025 80.925 ;
        RECT 78.085 80.665 78.345 80.925 ;
        RECT 78.620 80.715 78.880 80.975 ;
        RECT 75.795 80.235 76.055 80.495 ;
        RECT 76.115 80.235 76.375 80.495 ;
        RECT 76.435 80.235 76.695 80.495 ;
        RECT 77.530 80.235 77.790 80.495 ;
        RECT 77.850 80.235 78.110 80.495 ;
        RECT 78.620 80.395 78.880 80.655 ;
        RECT 72.495 79.805 72.755 80.065 ;
        RECT 72.815 79.805 73.075 80.065 ;
        RECT 73.135 79.805 73.395 80.065 ;
        RECT 78.620 80.075 78.880 80.335 ;
        RECT 75.795 79.805 76.055 80.065 ;
        RECT 76.115 79.805 76.375 80.065 ;
        RECT 76.435 79.805 76.695 80.065 ;
        RECT 77.445 79.805 77.705 80.065 ;
        RECT 77.765 79.805 78.025 80.065 ;
        RECT 78.085 79.805 78.345 80.065 ;
        RECT 78.620 79.755 78.880 80.015 ;
        RECT 72.730 79.375 72.990 79.635 ;
        RECT 73.050 79.375 73.310 79.635 ;
        RECT 75.795 79.375 76.055 79.635 ;
        RECT 76.115 79.375 76.375 79.635 ;
        RECT 76.435 79.375 76.695 79.635 ;
        RECT 77.530 79.375 77.790 79.635 ;
        RECT 77.850 79.375 78.110 79.635 ;
        RECT 72.730 78.945 72.990 79.205 ;
        RECT 73.050 78.945 73.310 79.205 ;
        RECT 72.730 78.515 72.990 78.775 ;
        RECT 73.050 78.515 73.310 78.775 ;
        RECT 72.730 77.865 72.990 78.125 ;
        RECT 73.050 77.865 73.310 78.125 ;
        RECT 75.955 78.945 76.215 79.205 ;
        RECT 76.275 78.945 76.535 79.205 ;
        RECT 77.530 78.945 77.790 79.205 ;
        RECT 77.850 78.945 78.110 79.205 ;
        RECT 75.955 78.515 76.215 78.775 ;
        RECT 76.275 78.515 76.535 78.775 ;
        RECT 77.530 78.515 77.790 78.775 ;
        RECT 77.850 78.515 78.110 78.775 ;
        RECT 75.955 77.865 76.215 78.125 ;
        RECT 76.275 77.865 76.535 78.125 ;
        RECT 77.530 77.865 77.790 78.125 ;
        RECT 77.850 77.865 78.110 78.125 ;
        RECT 80.450 81.955 80.710 82.215 ;
        RECT 80.770 81.955 81.030 82.215 ;
        RECT 82.025 81.955 82.285 82.215 ;
        RECT 82.345 81.955 82.605 82.215 ;
        RECT 80.450 81.525 80.710 81.785 ;
        RECT 80.770 81.525 81.030 81.785 ;
        RECT 82.025 81.525 82.285 81.785 ;
        RECT 82.345 81.525 82.605 81.785 ;
        RECT 83.835 81.745 84.095 82.005 ;
        RECT 83.835 81.425 84.095 81.685 ;
        RECT 80.450 81.095 80.710 81.355 ;
        RECT 80.770 81.095 81.030 81.355 ;
        RECT 81.865 81.095 82.125 81.355 ;
        RECT 82.185 81.095 82.445 81.355 ;
        RECT 82.505 81.095 82.765 81.355 ;
        RECT 79.680 80.715 79.940 80.975 ;
        RECT 80.215 80.665 80.475 80.925 ;
        RECT 80.535 80.665 80.795 80.925 ;
        RECT 80.855 80.665 81.115 80.925 ;
        RECT 81.865 80.665 82.125 80.925 ;
        RECT 82.185 80.665 82.445 80.925 ;
        RECT 82.505 80.665 82.765 80.925 ;
        RECT 79.680 80.395 79.940 80.655 ;
        RECT 79.680 80.075 79.940 80.335 ;
        RECT 80.450 80.235 80.710 80.495 ;
        RECT 80.770 80.235 81.030 80.495 ;
        RECT 81.865 80.235 82.125 80.495 ;
        RECT 82.185 80.235 82.445 80.495 ;
        RECT 82.505 80.235 82.765 80.495 ;
        RECT 85.250 81.955 85.510 82.215 ;
        RECT 85.570 81.955 85.830 82.215 ;
        RECT 85.250 81.525 85.510 81.785 ;
        RECT 85.570 81.525 85.830 81.785 ;
        RECT 85.250 81.095 85.510 81.355 ;
        RECT 85.570 81.095 85.830 81.355 ;
        RECT 85.165 80.665 85.425 80.925 ;
        RECT 85.485 80.665 85.745 80.925 ;
        RECT 85.805 80.665 86.065 80.925 ;
        RECT 86.340 80.825 86.600 81.085 ;
        RECT 86.340 80.505 86.600 80.765 ;
        RECT 85.250 80.235 85.510 80.495 ;
        RECT 85.570 80.235 85.830 80.495 ;
        RECT 79.680 79.755 79.940 80.015 ;
        RECT 80.215 79.805 80.475 80.065 ;
        RECT 80.535 79.805 80.795 80.065 ;
        RECT 80.855 79.805 81.115 80.065 ;
        RECT 81.865 79.805 82.125 80.065 ;
        RECT 82.185 79.805 82.445 80.065 ;
        RECT 82.505 79.805 82.765 80.065 ;
        RECT 85.165 79.805 85.425 80.065 ;
        RECT 85.485 79.805 85.745 80.065 ;
        RECT 85.805 79.805 86.065 80.065 ;
        RECT 80.450 79.375 80.710 79.635 ;
        RECT 80.770 79.375 81.030 79.635 ;
        RECT 81.865 79.375 82.125 79.635 ;
        RECT 82.185 79.375 82.445 79.635 ;
        RECT 82.505 79.375 82.765 79.635 ;
        RECT 85.250 79.375 85.510 79.635 ;
        RECT 85.570 79.375 85.830 79.635 ;
        RECT 80.450 78.945 80.710 79.205 ;
        RECT 80.770 78.945 81.030 79.205 ;
        RECT 82.025 78.945 82.285 79.205 ;
        RECT 82.345 78.945 82.605 79.205 ;
        RECT 80.450 78.515 80.710 78.775 ;
        RECT 80.770 78.515 81.030 78.775 ;
        RECT 82.025 78.515 82.285 78.775 ;
        RECT 82.345 78.515 82.605 78.775 ;
        RECT 80.450 77.865 80.710 78.125 ;
        RECT 80.770 77.865 81.030 78.125 ;
        RECT 82.025 77.865 82.285 78.125 ;
        RECT 82.345 77.865 82.605 78.125 ;
        RECT 85.250 78.945 85.510 79.205 ;
        RECT 85.570 78.945 85.830 79.205 ;
        RECT 85.250 78.515 85.510 78.775 ;
        RECT 85.570 78.515 85.830 78.775 ;
        RECT 85.250 77.865 85.510 78.125 ;
        RECT 85.570 77.865 85.830 78.125 ;
        RECT 89.160 82.305 89.420 82.565 ;
        RECT 89.480 82.305 89.740 82.565 ;
        RECT 89.800 82.305 90.060 82.565 ;
        RECT 89.160 81.875 89.420 82.135 ;
        RECT 89.480 81.875 89.740 82.135 ;
        RECT 89.800 81.875 90.060 82.135 ;
        RECT 91.155 82.210 91.415 82.470 ;
        RECT 91.155 81.890 91.415 82.150 ;
        RECT 89.160 81.445 89.420 81.705 ;
        RECT 89.480 81.445 89.740 81.705 ;
        RECT 89.800 81.445 90.060 81.705 ;
        RECT 89.160 81.015 89.420 81.275 ;
        RECT 89.480 81.015 89.740 81.275 ;
        RECT 89.800 81.015 90.060 81.275 ;
        RECT 93.010 82.305 93.270 82.565 ;
        RECT 93.330 82.305 93.590 82.565 ;
        RECT 93.650 82.305 93.910 82.565 ;
        RECT 93.010 81.875 93.270 82.135 ;
        RECT 93.330 81.875 93.590 82.135 ;
        RECT 93.650 81.875 93.910 82.135 ;
        RECT 93.010 81.445 93.270 81.705 ;
        RECT 93.330 81.445 93.590 81.705 ;
        RECT 93.650 81.445 93.910 81.705 ;
        RECT 92.530 81.015 92.790 81.275 ;
        RECT 92.850 81.015 93.110 81.275 ;
        RECT 93.170 81.015 93.430 81.275 ;
        RECT 93.490 81.015 93.750 81.275 ;
        RECT 93.810 81.015 94.070 81.275 ;
        RECT 94.130 81.015 94.390 81.275 ;
        RECT 89.160 80.585 89.420 80.845 ;
        RECT 89.480 80.585 89.740 80.845 ;
        RECT 89.800 80.585 90.060 80.845 ;
        RECT 93.010 80.585 93.270 80.845 ;
        RECT 93.330 80.585 93.590 80.845 ;
        RECT 93.650 80.585 93.910 80.845 ;
        RECT 89.160 80.155 89.420 80.415 ;
        RECT 89.480 80.155 89.740 80.415 ;
        RECT 89.800 80.155 90.060 80.415 ;
        RECT 92.530 80.155 92.790 80.415 ;
        RECT 92.850 80.155 93.110 80.415 ;
        RECT 93.170 80.155 93.430 80.415 ;
        RECT 93.490 80.155 93.750 80.415 ;
        RECT 93.810 80.155 94.070 80.415 ;
        RECT 94.130 80.155 94.390 80.415 ;
        RECT 89.160 79.725 89.420 79.985 ;
        RECT 89.480 79.725 89.740 79.985 ;
        RECT 89.800 79.725 90.060 79.985 ;
        RECT 93.010 79.725 93.270 79.985 ;
        RECT 93.330 79.725 93.590 79.985 ;
        RECT 93.650 79.725 93.910 79.985 ;
        RECT 89.160 79.295 89.420 79.555 ;
        RECT 89.480 79.295 89.740 79.555 ;
        RECT 89.800 79.295 90.060 79.555 ;
        RECT 89.160 78.865 89.420 79.125 ;
        RECT 89.480 78.865 89.740 79.125 ;
        RECT 89.800 78.865 90.060 79.125 ;
        RECT 93.010 79.295 93.270 79.555 ;
        RECT 93.330 79.295 93.590 79.555 ;
        RECT 93.650 79.295 93.910 79.555 ;
        RECT 93.010 78.865 93.270 79.125 ;
        RECT 93.330 78.865 93.590 79.125 ;
        RECT 93.650 78.865 93.910 79.125 ;
        RECT 89.160 78.195 89.420 78.455 ;
        RECT 89.480 78.195 89.740 78.455 ;
        RECT 89.800 78.195 90.060 78.455 ;
        RECT 93.010 78.195 93.270 78.455 ;
        RECT 93.330 78.195 93.590 78.455 ;
        RECT 93.650 78.195 93.910 78.455 ;
        RECT 65.380 72.315 65.640 72.575 ;
        RECT 65.700 72.315 65.960 72.575 ;
        RECT 66.020 72.315 66.280 72.575 ;
        RECT 69.230 72.315 69.490 72.575 ;
        RECT 69.550 72.315 69.810 72.575 ;
        RECT 69.870 72.315 70.130 72.575 ;
        RECT 65.380 71.645 65.640 71.905 ;
        RECT 65.700 71.645 65.960 71.905 ;
        RECT 66.020 71.645 66.280 71.905 ;
        RECT 65.380 71.215 65.640 71.475 ;
        RECT 65.700 71.215 65.960 71.475 ;
        RECT 66.020 71.215 66.280 71.475 ;
        RECT 67.375 71.550 67.635 71.810 ;
        RECT 67.375 71.230 67.635 71.490 ;
        RECT 65.380 70.785 65.640 71.045 ;
        RECT 65.700 70.785 65.960 71.045 ;
        RECT 66.020 70.785 66.280 71.045 ;
        RECT 65.380 70.355 65.640 70.615 ;
        RECT 65.700 70.355 65.960 70.615 ;
        RECT 66.020 70.355 66.280 70.615 ;
        RECT 69.230 71.645 69.490 71.905 ;
        RECT 69.550 71.645 69.810 71.905 ;
        RECT 69.870 71.645 70.130 71.905 ;
        RECT 69.230 71.215 69.490 71.475 ;
        RECT 69.550 71.215 69.810 71.475 ;
        RECT 69.870 71.215 70.130 71.475 ;
        RECT 69.230 70.785 69.490 71.045 ;
        RECT 69.550 70.785 69.810 71.045 ;
        RECT 69.870 70.785 70.130 71.045 ;
        RECT 68.750 70.355 69.010 70.615 ;
        RECT 69.070 70.355 69.330 70.615 ;
        RECT 69.390 70.355 69.650 70.615 ;
        RECT 69.710 70.355 69.970 70.615 ;
        RECT 70.030 70.355 70.290 70.615 ;
        RECT 70.350 70.355 70.610 70.615 ;
        RECT 65.380 69.925 65.640 70.185 ;
        RECT 65.700 69.925 65.960 70.185 ;
        RECT 66.020 69.925 66.280 70.185 ;
        RECT 69.230 69.925 69.490 70.185 ;
        RECT 69.550 69.925 69.810 70.185 ;
        RECT 69.870 69.925 70.130 70.185 ;
        RECT 65.380 69.495 65.640 69.755 ;
        RECT 65.700 69.495 65.960 69.755 ;
        RECT 66.020 69.495 66.280 69.755 ;
        RECT 67.055 69.495 67.315 69.755 ;
        RECT 67.375 69.495 67.635 69.755 ;
        RECT 67.695 69.495 67.955 69.755 ;
        RECT 65.380 69.065 65.640 69.325 ;
        RECT 65.700 69.065 65.960 69.325 ;
        RECT 66.020 69.065 66.280 69.325 ;
        RECT 65.380 68.635 65.640 68.895 ;
        RECT 65.700 68.635 65.960 68.895 ;
        RECT 66.020 68.635 66.280 68.895 ;
        RECT 65.380 68.205 65.640 68.465 ;
        RECT 65.700 68.205 65.960 68.465 ;
        RECT 66.020 68.205 66.280 68.465 ;
        RECT 65.380 67.775 65.640 68.035 ;
        RECT 65.700 67.775 65.960 68.035 ;
        RECT 66.020 67.775 66.280 68.035 ;
        RECT 65.380 67.345 65.640 67.605 ;
        RECT 65.700 67.345 65.960 67.605 ;
        RECT 66.020 67.345 66.280 67.605 ;
        RECT 68.750 69.495 69.010 69.755 ;
        RECT 69.070 69.495 69.330 69.755 ;
        RECT 69.390 69.495 69.650 69.755 ;
        RECT 69.710 69.495 69.970 69.755 ;
        RECT 70.030 69.495 70.290 69.755 ;
        RECT 70.350 69.495 70.610 69.755 ;
        RECT 69.230 69.065 69.490 69.325 ;
        RECT 69.550 69.065 69.810 69.325 ;
        RECT 69.870 69.065 70.130 69.325 ;
        RECT 68.750 68.635 69.010 68.895 ;
        RECT 69.070 68.635 69.330 68.895 ;
        RECT 69.390 68.635 69.650 68.895 ;
        RECT 69.710 68.635 69.970 68.895 ;
        RECT 70.030 68.635 70.290 68.895 ;
        RECT 70.350 68.635 70.610 68.895 ;
        RECT 69.230 68.205 69.490 68.465 ;
        RECT 69.550 68.205 69.810 68.465 ;
        RECT 69.870 68.205 70.130 68.465 ;
        RECT 68.750 67.775 69.010 68.035 ;
        RECT 69.070 67.775 69.330 68.035 ;
        RECT 69.390 67.775 69.650 68.035 ;
        RECT 69.710 67.775 69.970 68.035 ;
        RECT 70.030 67.775 70.290 68.035 ;
        RECT 70.350 67.775 70.610 68.035 ;
        RECT 69.230 67.345 69.490 67.605 ;
        RECT 69.550 67.345 69.810 67.605 ;
        RECT 69.870 67.345 70.130 67.605 ;
        RECT 65.380 66.915 65.640 67.175 ;
        RECT 65.700 66.915 65.960 67.175 ;
        RECT 66.020 66.915 66.280 67.175 ;
        RECT 68.750 66.915 69.010 67.175 ;
        RECT 69.070 66.915 69.330 67.175 ;
        RECT 69.390 66.915 69.650 67.175 ;
        RECT 69.710 66.915 69.970 67.175 ;
        RECT 70.030 66.915 70.290 67.175 ;
        RECT 70.350 66.915 70.610 67.175 ;
        RECT 65.380 66.485 65.640 66.745 ;
        RECT 65.700 66.485 65.960 66.745 ;
        RECT 66.020 66.485 66.280 66.745 ;
        RECT 65.380 66.055 65.640 66.315 ;
        RECT 65.700 66.055 65.960 66.315 ;
        RECT 66.020 66.055 66.280 66.315 ;
        RECT 65.380 65.625 65.640 65.885 ;
        RECT 65.700 65.625 65.960 65.885 ;
        RECT 66.020 65.625 66.280 65.885 ;
        RECT 65.380 65.195 65.640 65.455 ;
        RECT 65.700 65.195 65.960 65.455 ;
        RECT 66.020 65.195 66.280 65.455 ;
        RECT 69.230 66.485 69.490 66.745 ;
        RECT 69.550 66.485 69.810 66.745 ;
        RECT 69.870 66.485 70.130 66.745 ;
        RECT 68.750 66.055 69.010 66.315 ;
        RECT 69.070 66.055 69.330 66.315 ;
        RECT 69.390 66.055 69.650 66.315 ;
        RECT 69.710 66.055 69.970 66.315 ;
        RECT 70.030 66.055 70.290 66.315 ;
        RECT 70.350 66.055 70.610 66.315 ;
        RECT 69.230 65.625 69.490 65.885 ;
        RECT 69.550 65.625 69.810 65.885 ;
        RECT 69.870 65.625 70.130 65.885 ;
        RECT 68.750 65.195 69.010 65.455 ;
        RECT 69.070 65.195 69.330 65.455 ;
        RECT 69.390 65.195 69.650 65.455 ;
        RECT 69.710 65.195 69.970 65.455 ;
        RECT 70.030 65.195 70.290 65.455 ;
        RECT 70.350 65.195 70.610 65.455 ;
        RECT 65.380 64.765 65.640 65.025 ;
        RECT 65.700 64.765 65.960 65.025 ;
        RECT 66.020 64.765 66.280 65.025 ;
        RECT 69.230 64.765 69.490 65.025 ;
        RECT 69.550 64.765 69.810 65.025 ;
        RECT 69.870 64.765 70.130 65.025 ;
        RECT 65.380 64.335 65.640 64.595 ;
        RECT 65.700 64.335 65.960 64.595 ;
        RECT 66.020 64.335 66.280 64.595 ;
        RECT 65.380 63.905 65.640 64.165 ;
        RECT 65.700 63.905 65.960 64.165 ;
        RECT 66.020 63.905 66.280 64.165 ;
        RECT 69.230 64.335 69.490 64.595 ;
        RECT 69.550 64.335 69.810 64.595 ;
        RECT 69.870 64.335 70.130 64.595 ;
        RECT 69.230 63.905 69.490 64.165 ;
        RECT 69.550 63.905 69.810 64.165 ;
        RECT 69.870 63.905 70.130 64.165 ;
        RECT 65.380 63.235 65.640 63.495 ;
        RECT 65.700 63.235 65.960 63.495 ;
        RECT 66.020 63.235 66.280 63.495 ;
        RECT 69.230 63.235 69.490 63.495 ;
        RECT 69.550 63.235 69.810 63.495 ;
        RECT 69.870 63.235 70.130 63.495 ;
        RECT 74.400 72.315 74.660 72.575 ;
        RECT 74.720 72.315 74.980 72.575 ;
        RECT 75.040 72.315 75.300 72.575 ;
        RECT 78.250 72.315 78.510 72.575 ;
        RECT 78.570 72.315 78.830 72.575 ;
        RECT 78.890 72.315 79.150 72.575 ;
        RECT 81.340 72.315 81.600 72.575 ;
        RECT 81.660 72.315 81.920 72.575 ;
        RECT 81.980 72.315 82.240 72.575 ;
        RECT 85.190 72.315 85.450 72.575 ;
        RECT 85.510 72.315 85.770 72.575 ;
        RECT 85.830 72.315 86.090 72.575 ;
        RECT 74.400 71.645 74.660 71.905 ;
        RECT 74.720 71.645 74.980 71.905 ;
        RECT 75.040 71.645 75.300 71.905 ;
        RECT 74.400 71.215 74.660 71.475 ;
        RECT 74.720 71.215 74.980 71.475 ;
        RECT 75.040 71.215 75.300 71.475 ;
        RECT 76.395 71.550 76.655 71.810 ;
        RECT 76.395 71.230 76.655 71.490 ;
        RECT 74.400 70.785 74.660 71.045 ;
        RECT 74.720 70.785 74.980 71.045 ;
        RECT 75.040 70.785 75.300 71.045 ;
        RECT 74.400 70.355 74.660 70.615 ;
        RECT 74.720 70.355 74.980 70.615 ;
        RECT 75.040 70.355 75.300 70.615 ;
        RECT 78.250 71.645 78.510 71.905 ;
        RECT 78.570 71.645 78.830 71.905 ;
        RECT 78.890 71.645 79.150 71.905 ;
        RECT 78.250 71.215 78.510 71.475 ;
        RECT 78.570 71.215 78.830 71.475 ;
        RECT 78.890 71.215 79.150 71.475 ;
        RECT 78.250 70.785 78.510 71.045 ;
        RECT 78.570 70.785 78.830 71.045 ;
        RECT 78.890 70.785 79.150 71.045 ;
        RECT 77.770 70.355 78.030 70.615 ;
        RECT 78.090 70.355 78.350 70.615 ;
        RECT 78.410 70.355 78.670 70.615 ;
        RECT 78.730 70.355 78.990 70.615 ;
        RECT 79.050 70.355 79.310 70.615 ;
        RECT 79.370 70.355 79.630 70.615 ;
        RECT 74.400 69.925 74.660 70.185 ;
        RECT 74.720 69.925 74.980 70.185 ;
        RECT 75.040 69.925 75.300 70.185 ;
        RECT 78.250 69.925 78.510 70.185 ;
        RECT 78.570 69.925 78.830 70.185 ;
        RECT 78.890 69.925 79.150 70.185 ;
        RECT 74.400 69.495 74.660 69.755 ;
        RECT 74.720 69.495 74.980 69.755 ;
        RECT 75.040 69.495 75.300 69.755 ;
        RECT 76.075 69.495 76.335 69.755 ;
        RECT 76.395 69.495 76.655 69.755 ;
        RECT 76.715 69.495 76.975 69.755 ;
        RECT 74.400 69.065 74.660 69.325 ;
        RECT 74.720 69.065 74.980 69.325 ;
        RECT 75.040 69.065 75.300 69.325 ;
        RECT 74.400 68.635 74.660 68.895 ;
        RECT 74.720 68.635 74.980 68.895 ;
        RECT 75.040 68.635 75.300 68.895 ;
        RECT 74.400 68.205 74.660 68.465 ;
        RECT 74.720 68.205 74.980 68.465 ;
        RECT 75.040 68.205 75.300 68.465 ;
        RECT 74.400 67.775 74.660 68.035 ;
        RECT 74.720 67.775 74.980 68.035 ;
        RECT 75.040 67.775 75.300 68.035 ;
        RECT 74.400 67.345 74.660 67.605 ;
        RECT 74.720 67.345 74.980 67.605 ;
        RECT 75.040 67.345 75.300 67.605 ;
        RECT 77.770 69.495 78.030 69.755 ;
        RECT 78.090 69.495 78.350 69.755 ;
        RECT 78.410 69.495 78.670 69.755 ;
        RECT 78.730 69.495 78.990 69.755 ;
        RECT 79.050 69.495 79.310 69.755 ;
        RECT 79.370 69.495 79.630 69.755 ;
        RECT 78.250 69.065 78.510 69.325 ;
        RECT 78.570 69.065 78.830 69.325 ;
        RECT 78.890 69.065 79.150 69.325 ;
        RECT 77.770 68.635 78.030 68.895 ;
        RECT 78.090 68.635 78.350 68.895 ;
        RECT 78.410 68.635 78.670 68.895 ;
        RECT 78.730 68.635 78.990 68.895 ;
        RECT 79.050 68.635 79.310 68.895 ;
        RECT 79.370 68.635 79.630 68.895 ;
        RECT 78.250 68.205 78.510 68.465 ;
        RECT 78.570 68.205 78.830 68.465 ;
        RECT 78.890 68.205 79.150 68.465 ;
        RECT 77.770 67.775 78.030 68.035 ;
        RECT 78.090 67.775 78.350 68.035 ;
        RECT 78.410 67.775 78.670 68.035 ;
        RECT 78.730 67.775 78.990 68.035 ;
        RECT 79.050 67.775 79.310 68.035 ;
        RECT 79.370 67.775 79.630 68.035 ;
        RECT 78.250 67.345 78.510 67.605 ;
        RECT 78.570 67.345 78.830 67.605 ;
        RECT 78.890 67.345 79.150 67.605 ;
        RECT 74.400 66.915 74.660 67.175 ;
        RECT 74.720 66.915 74.980 67.175 ;
        RECT 75.040 66.915 75.300 67.175 ;
        RECT 77.770 66.915 78.030 67.175 ;
        RECT 78.090 66.915 78.350 67.175 ;
        RECT 78.410 66.915 78.670 67.175 ;
        RECT 78.730 66.915 78.990 67.175 ;
        RECT 79.050 66.915 79.310 67.175 ;
        RECT 79.370 66.915 79.630 67.175 ;
        RECT 74.400 66.485 74.660 66.745 ;
        RECT 74.720 66.485 74.980 66.745 ;
        RECT 75.040 66.485 75.300 66.745 ;
        RECT 74.400 66.055 74.660 66.315 ;
        RECT 74.720 66.055 74.980 66.315 ;
        RECT 75.040 66.055 75.300 66.315 ;
        RECT 74.400 65.625 74.660 65.885 ;
        RECT 74.720 65.625 74.980 65.885 ;
        RECT 75.040 65.625 75.300 65.885 ;
        RECT 74.400 65.195 74.660 65.455 ;
        RECT 74.720 65.195 74.980 65.455 ;
        RECT 75.040 65.195 75.300 65.455 ;
        RECT 78.250 66.485 78.510 66.745 ;
        RECT 78.570 66.485 78.830 66.745 ;
        RECT 78.890 66.485 79.150 66.745 ;
        RECT 77.770 66.055 78.030 66.315 ;
        RECT 78.090 66.055 78.350 66.315 ;
        RECT 78.410 66.055 78.670 66.315 ;
        RECT 78.730 66.055 78.990 66.315 ;
        RECT 79.050 66.055 79.310 66.315 ;
        RECT 79.370 66.055 79.630 66.315 ;
        RECT 78.250 65.625 78.510 65.885 ;
        RECT 78.570 65.625 78.830 65.885 ;
        RECT 78.890 65.625 79.150 65.885 ;
        RECT 77.770 65.195 78.030 65.455 ;
        RECT 78.090 65.195 78.350 65.455 ;
        RECT 78.410 65.195 78.670 65.455 ;
        RECT 78.730 65.195 78.990 65.455 ;
        RECT 79.050 65.195 79.310 65.455 ;
        RECT 79.370 65.195 79.630 65.455 ;
        RECT 74.400 64.765 74.660 65.025 ;
        RECT 74.720 64.765 74.980 65.025 ;
        RECT 75.040 64.765 75.300 65.025 ;
        RECT 78.250 64.765 78.510 65.025 ;
        RECT 78.570 64.765 78.830 65.025 ;
        RECT 78.890 64.765 79.150 65.025 ;
        RECT 74.400 64.335 74.660 64.595 ;
        RECT 74.720 64.335 74.980 64.595 ;
        RECT 75.040 64.335 75.300 64.595 ;
        RECT 74.400 63.905 74.660 64.165 ;
        RECT 74.720 63.905 74.980 64.165 ;
        RECT 75.040 63.905 75.300 64.165 ;
        RECT 78.250 64.335 78.510 64.595 ;
        RECT 78.570 64.335 78.830 64.595 ;
        RECT 78.890 64.335 79.150 64.595 ;
        RECT 78.250 63.905 78.510 64.165 ;
        RECT 78.570 63.905 78.830 64.165 ;
        RECT 78.890 63.905 79.150 64.165 ;
        RECT 81.340 71.645 81.600 71.905 ;
        RECT 81.660 71.645 81.920 71.905 ;
        RECT 81.980 71.645 82.240 71.905 ;
        RECT 81.340 71.215 81.600 71.475 ;
        RECT 81.660 71.215 81.920 71.475 ;
        RECT 81.980 71.215 82.240 71.475 ;
        RECT 83.835 71.550 84.095 71.810 ;
        RECT 83.835 71.230 84.095 71.490 ;
        RECT 81.340 70.785 81.600 71.045 ;
        RECT 81.660 70.785 81.920 71.045 ;
        RECT 81.980 70.785 82.240 71.045 ;
        RECT 80.860 70.355 81.120 70.615 ;
        RECT 81.180 70.355 81.440 70.615 ;
        RECT 81.500 70.355 81.760 70.615 ;
        RECT 81.820 70.355 82.080 70.615 ;
        RECT 82.140 70.355 82.400 70.615 ;
        RECT 82.460 70.355 82.720 70.615 ;
        RECT 85.190 71.645 85.450 71.905 ;
        RECT 85.510 71.645 85.770 71.905 ;
        RECT 85.830 71.645 86.090 71.905 ;
        RECT 85.190 71.215 85.450 71.475 ;
        RECT 85.510 71.215 85.770 71.475 ;
        RECT 85.830 71.215 86.090 71.475 ;
        RECT 85.190 70.785 85.450 71.045 ;
        RECT 85.510 70.785 85.770 71.045 ;
        RECT 85.830 70.785 86.090 71.045 ;
        RECT 85.190 70.355 85.450 70.615 ;
        RECT 85.510 70.355 85.770 70.615 ;
        RECT 85.830 70.355 86.090 70.615 ;
        RECT 81.340 69.925 81.600 70.185 ;
        RECT 81.660 69.925 81.920 70.185 ;
        RECT 81.980 69.925 82.240 70.185 ;
        RECT 85.190 69.925 85.450 70.185 ;
        RECT 85.510 69.925 85.770 70.185 ;
        RECT 85.830 69.925 86.090 70.185 ;
        RECT 80.860 69.495 81.120 69.755 ;
        RECT 81.180 69.495 81.440 69.755 ;
        RECT 81.500 69.495 81.760 69.755 ;
        RECT 81.820 69.495 82.080 69.755 ;
        RECT 82.140 69.495 82.400 69.755 ;
        RECT 82.460 69.495 82.720 69.755 ;
        RECT 83.515 69.495 83.775 69.755 ;
        RECT 83.835 69.495 84.095 69.755 ;
        RECT 84.155 69.495 84.415 69.755 ;
        RECT 81.340 69.065 81.600 69.325 ;
        RECT 81.660 69.065 81.920 69.325 ;
        RECT 81.980 69.065 82.240 69.325 ;
        RECT 80.860 68.635 81.120 68.895 ;
        RECT 81.180 68.635 81.440 68.895 ;
        RECT 81.500 68.635 81.760 68.895 ;
        RECT 81.820 68.635 82.080 68.895 ;
        RECT 82.140 68.635 82.400 68.895 ;
        RECT 82.460 68.635 82.720 68.895 ;
        RECT 81.340 68.205 81.600 68.465 ;
        RECT 81.660 68.205 81.920 68.465 ;
        RECT 81.980 68.205 82.240 68.465 ;
        RECT 80.860 67.775 81.120 68.035 ;
        RECT 81.180 67.775 81.440 68.035 ;
        RECT 81.500 67.775 81.760 68.035 ;
        RECT 81.820 67.775 82.080 68.035 ;
        RECT 82.140 67.775 82.400 68.035 ;
        RECT 82.460 67.775 82.720 68.035 ;
        RECT 81.340 67.345 81.600 67.605 ;
        RECT 81.660 67.345 81.920 67.605 ;
        RECT 81.980 67.345 82.240 67.605 ;
        RECT 85.190 69.495 85.450 69.755 ;
        RECT 85.510 69.495 85.770 69.755 ;
        RECT 85.830 69.495 86.090 69.755 ;
        RECT 85.190 69.065 85.450 69.325 ;
        RECT 85.510 69.065 85.770 69.325 ;
        RECT 85.830 69.065 86.090 69.325 ;
        RECT 85.190 68.635 85.450 68.895 ;
        RECT 85.510 68.635 85.770 68.895 ;
        RECT 85.830 68.635 86.090 68.895 ;
        RECT 85.190 68.205 85.450 68.465 ;
        RECT 85.510 68.205 85.770 68.465 ;
        RECT 85.830 68.205 86.090 68.465 ;
        RECT 85.190 67.775 85.450 68.035 ;
        RECT 85.510 67.775 85.770 68.035 ;
        RECT 85.830 67.775 86.090 68.035 ;
        RECT 85.190 67.345 85.450 67.605 ;
        RECT 85.510 67.345 85.770 67.605 ;
        RECT 85.830 67.345 86.090 67.605 ;
        RECT 80.860 66.915 81.120 67.175 ;
        RECT 81.180 66.915 81.440 67.175 ;
        RECT 81.500 66.915 81.760 67.175 ;
        RECT 81.820 66.915 82.080 67.175 ;
        RECT 82.140 66.915 82.400 67.175 ;
        RECT 82.460 66.915 82.720 67.175 ;
        RECT 85.190 66.915 85.450 67.175 ;
        RECT 85.510 66.915 85.770 67.175 ;
        RECT 85.830 66.915 86.090 67.175 ;
        RECT 81.340 66.485 81.600 66.745 ;
        RECT 81.660 66.485 81.920 66.745 ;
        RECT 81.980 66.485 82.240 66.745 ;
        RECT 80.860 66.055 81.120 66.315 ;
        RECT 81.180 66.055 81.440 66.315 ;
        RECT 81.500 66.055 81.760 66.315 ;
        RECT 81.820 66.055 82.080 66.315 ;
        RECT 82.140 66.055 82.400 66.315 ;
        RECT 82.460 66.055 82.720 66.315 ;
        RECT 81.340 65.625 81.600 65.885 ;
        RECT 81.660 65.625 81.920 65.885 ;
        RECT 81.980 65.625 82.240 65.885 ;
        RECT 80.860 65.195 81.120 65.455 ;
        RECT 81.180 65.195 81.440 65.455 ;
        RECT 81.500 65.195 81.760 65.455 ;
        RECT 81.820 65.195 82.080 65.455 ;
        RECT 82.140 65.195 82.400 65.455 ;
        RECT 82.460 65.195 82.720 65.455 ;
        RECT 85.190 66.485 85.450 66.745 ;
        RECT 85.510 66.485 85.770 66.745 ;
        RECT 85.830 66.485 86.090 66.745 ;
        RECT 85.190 66.055 85.450 66.315 ;
        RECT 85.510 66.055 85.770 66.315 ;
        RECT 85.830 66.055 86.090 66.315 ;
        RECT 85.190 65.625 85.450 65.885 ;
        RECT 85.510 65.625 85.770 65.885 ;
        RECT 85.830 65.625 86.090 65.885 ;
        RECT 85.190 65.195 85.450 65.455 ;
        RECT 85.510 65.195 85.770 65.455 ;
        RECT 85.830 65.195 86.090 65.455 ;
        RECT 81.340 64.765 81.600 65.025 ;
        RECT 81.660 64.765 81.920 65.025 ;
        RECT 81.980 64.765 82.240 65.025 ;
        RECT 85.190 64.765 85.450 65.025 ;
        RECT 85.510 64.765 85.770 65.025 ;
        RECT 85.830 64.765 86.090 65.025 ;
        RECT 81.340 64.335 81.600 64.595 ;
        RECT 81.660 64.335 81.920 64.595 ;
        RECT 81.980 64.335 82.240 64.595 ;
        RECT 81.340 63.905 81.600 64.165 ;
        RECT 81.660 63.905 81.920 64.165 ;
        RECT 81.980 63.905 82.240 64.165 ;
        RECT 85.190 64.335 85.450 64.595 ;
        RECT 85.510 64.335 85.770 64.595 ;
        RECT 85.830 64.335 86.090 64.595 ;
        RECT 85.190 63.905 85.450 64.165 ;
        RECT 85.510 63.905 85.770 64.165 ;
        RECT 85.830 63.905 86.090 64.165 ;
        RECT 74.400 63.235 74.660 63.495 ;
        RECT 74.720 63.235 74.980 63.495 ;
        RECT 75.040 63.235 75.300 63.495 ;
        RECT 78.250 63.235 78.510 63.495 ;
        RECT 78.570 63.235 78.830 63.495 ;
        RECT 78.890 63.235 79.150 63.495 ;
        RECT 81.340 63.235 81.600 63.495 ;
        RECT 81.660 63.235 81.920 63.495 ;
        RECT 81.980 63.235 82.240 63.495 ;
        RECT 85.190 63.235 85.450 63.495 ;
        RECT 85.510 63.235 85.770 63.495 ;
        RECT 85.830 63.235 86.090 63.495 ;
        RECT 89.160 72.315 89.420 72.575 ;
        RECT 89.480 72.315 89.740 72.575 ;
        RECT 89.800 72.315 90.060 72.575 ;
        RECT 93.010 72.315 93.270 72.575 ;
        RECT 93.330 72.315 93.590 72.575 ;
        RECT 93.650 72.315 93.910 72.575 ;
        RECT 89.160 71.645 89.420 71.905 ;
        RECT 89.480 71.645 89.740 71.905 ;
        RECT 89.800 71.645 90.060 71.905 ;
        RECT 89.160 71.215 89.420 71.475 ;
        RECT 89.480 71.215 89.740 71.475 ;
        RECT 89.800 71.215 90.060 71.475 ;
        RECT 91.155 71.550 91.415 71.810 ;
        RECT 91.155 71.230 91.415 71.490 ;
        RECT 89.160 70.785 89.420 71.045 ;
        RECT 89.480 70.785 89.740 71.045 ;
        RECT 89.800 70.785 90.060 71.045 ;
        RECT 89.160 70.355 89.420 70.615 ;
        RECT 89.480 70.355 89.740 70.615 ;
        RECT 89.800 70.355 90.060 70.615 ;
        RECT 93.010 71.645 93.270 71.905 ;
        RECT 93.330 71.645 93.590 71.905 ;
        RECT 93.650 71.645 93.910 71.905 ;
        RECT 93.010 71.215 93.270 71.475 ;
        RECT 93.330 71.215 93.590 71.475 ;
        RECT 93.650 71.215 93.910 71.475 ;
        RECT 93.010 70.785 93.270 71.045 ;
        RECT 93.330 70.785 93.590 71.045 ;
        RECT 93.650 70.785 93.910 71.045 ;
        RECT 92.530 70.355 92.790 70.615 ;
        RECT 92.850 70.355 93.110 70.615 ;
        RECT 93.170 70.355 93.430 70.615 ;
        RECT 93.490 70.355 93.750 70.615 ;
        RECT 93.810 70.355 94.070 70.615 ;
        RECT 94.130 70.355 94.390 70.615 ;
        RECT 89.160 69.925 89.420 70.185 ;
        RECT 89.480 69.925 89.740 70.185 ;
        RECT 89.800 69.925 90.060 70.185 ;
        RECT 93.010 69.925 93.270 70.185 ;
        RECT 93.330 69.925 93.590 70.185 ;
        RECT 93.650 69.925 93.910 70.185 ;
        RECT 89.160 69.495 89.420 69.755 ;
        RECT 89.480 69.495 89.740 69.755 ;
        RECT 89.800 69.495 90.060 69.755 ;
        RECT 90.835 69.495 91.095 69.755 ;
        RECT 91.155 69.495 91.415 69.755 ;
        RECT 91.475 69.495 91.735 69.755 ;
        RECT 89.160 69.065 89.420 69.325 ;
        RECT 89.480 69.065 89.740 69.325 ;
        RECT 89.800 69.065 90.060 69.325 ;
        RECT 89.160 68.635 89.420 68.895 ;
        RECT 89.480 68.635 89.740 68.895 ;
        RECT 89.800 68.635 90.060 68.895 ;
        RECT 89.160 68.205 89.420 68.465 ;
        RECT 89.480 68.205 89.740 68.465 ;
        RECT 89.800 68.205 90.060 68.465 ;
        RECT 89.160 67.775 89.420 68.035 ;
        RECT 89.480 67.775 89.740 68.035 ;
        RECT 89.800 67.775 90.060 68.035 ;
        RECT 89.160 67.345 89.420 67.605 ;
        RECT 89.480 67.345 89.740 67.605 ;
        RECT 89.800 67.345 90.060 67.605 ;
        RECT 92.530 69.495 92.790 69.755 ;
        RECT 92.850 69.495 93.110 69.755 ;
        RECT 93.170 69.495 93.430 69.755 ;
        RECT 93.490 69.495 93.750 69.755 ;
        RECT 93.810 69.495 94.070 69.755 ;
        RECT 94.130 69.495 94.390 69.755 ;
        RECT 93.010 69.065 93.270 69.325 ;
        RECT 93.330 69.065 93.590 69.325 ;
        RECT 93.650 69.065 93.910 69.325 ;
        RECT 92.530 68.635 92.790 68.895 ;
        RECT 92.850 68.635 93.110 68.895 ;
        RECT 93.170 68.635 93.430 68.895 ;
        RECT 93.490 68.635 93.750 68.895 ;
        RECT 93.810 68.635 94.070 68.895 ;
        RECT 94.130 68.635 94.390 68.895 ;
        RECT 93.010 68.205 93.270 68.465 ;
        RECT 93.330 68.205 93.590 68.465 ;
        RECT 93.650 68.205 93.910 68.465 ;
        RECT 92.530 67.775 92.790 68.035 ;
        RECT 92.850 67.775 93.110 68.035 ;
        RECT 93.170 67.775 93.430 68.035 ;
        RECT 93.490 67.775 93.750 68.035 ;
        RECT 93.810 67.775 94.070 68.035 ;
        RECT 94.130 67.775 94.390 68.035 ;
        RECT 93.010 67.345 93.270 67.605 ;
        RECT 93.330 67.345 93.590 67.605 ;
        RECT 93.650 67.345 93.910 67.605 ;
        RECT 89.160 66.915 89.420 67.175 ;
        RECT 89.480 66.915 89.740 67.175 ;
        RECT 89.800 66.915 90.060 67.175 ;
        RECT 92.530 66.915 92.790 67.175 ;
        RECT 92.850 66.915 93.110 67.175 ;
        RECT 93.170 66.915 93.430 67.175 ;
        RECT 93.490 66.915 93.750 67.175 ;
        RECT 93.810 66.915 94.070 67.175 ;
        RECT 94.130 66.915 94.390 67.175 ;
        RECT 89.160 66.485 89.420 66.745 ;
        RECT 89.480 66.485 89.740 66.745 ;
        RECT 89.800 66.485 90.060 66.745 ;
        RECT 89.160 66.055 89.420 66.315 ;
        RECT 89.480 66.055 89.740 66.315 ;
        RECT 89.800 66.055 90.060 66.315 ;
        RECT 89.160 65.625 89.420 65.885 ;
        RECT 89.480 65.625 89.740 65.885 ;
        RECT 89.800 65.625 90.060 65.885 ;
        RECT 89.160 65.195 89.420 65.455 ;
        RECT 89.480 65.195 89.740 65.455 ;
        RECT 89.800 65.195 90.060 65.455 ;
        RECT 93.010 66.485 93.270 66.745 ;
        RECT 93.330 66.485 93.590 66.745 ;
        RECT 93.650 66.485 93.910 66.745 ;
        RECT 92.530 66.055 92.790 66.315 ;
        RECT 92.850 66.055 93.110 66.315 ;
        RECT 93.170 66.055 93.430 66.315 ;
        RECT 93.490 66.055 93.750 66.315 ;
        RECT 93.810 66.055 94.070 66.315 ;
        RECT 94.130 66.055 94.390 66.315 ;
        RECT 93.010 65.625 93.270 65.885 ;
        RECT 93.330 65.625 93.590 65.885 ;
        RECT 93.650 65.625 93.910 65.885 ;
        RECT 92.530 65.195 92.790 65.455 ;
        RECT 92.850 65.195 93.110 65.455 ;
        RECT 93.170 65.195 93.430 65.455 ;
        RECT 93.490 65.195 93.750 65.455 ;
        RECT 93.810 65.195 94.070 65.455 ;
        RECT 94.130 65.195 94.390 65.455 ;
        RECT 89.160 64.765 89.420 65.025 ;
        RECT 89.480 64.765 89.740 65.025 ;
        RECT 89.800 64.765 90.060 65.025 ;
        RECT 93.010 64.765 93.270 65.025 ;
        RECT 93.330 64.765 93.590 65.025 ;
        RECT 93.650 64.765 93.910 65.025 ;
        RECT 89.160 64.335 89.420 64.595 ;
        RECT 89.480 64.335 89.740 64.595 ;
        RECT 89.800 64.335 90.060 64.595 ;
        RECT 89.160 63.905 89.420 64.165 ;
        RECT 89.480 63.905 89.740 64.165 ;
        RECT 89.800 63.905 90.060 64.165 ;
        RECT 93.010 64.335 93.270 64.595 ;
        RECT 93.330 64.335 93.590 64.595 ;
        RECT 93.650 64.335 93.910 64.595 ;
        RECT 93.010 63.905 93.270 64.165 ;
        RECT 93.330 63.905 93.590 64.165 ;
        RECT 93.650 63.905 93.910 64.165 ;
        RECT 89.160 63.235 89.420 63.495 ;
        RECT 89.480 63.235 89.740 63.495 ;
        RECT 89.800 63.235 90.060 63.495 ;
        RECT 93.010 63.235 93.270 63.495 ;
        RECT 93.330 63.235 93.590 63.495 ;
        RECT 93.650 63.235 93.910 63.495 ;
        RECT 109.665 164.035 109.925 164.295 ;
        RECT 109.985 164.035 110.245 164.295 ;
        RECT 109.665 161.755 109.925 162.015 ;
        RECT 109.985 161.755 110.245 162.015 ;
        RECT 111.035 164.035 111.295 164.295 ;
        RECT 111.355 164.035 111.615 164.295 ;
        RECT 111.035 161.755 111.295 162.015 ;
        RECT 111.355 161.755 111.615 162.015 ;
        RECT 112.405 164.035 112.665 164.295 ;
        RECT 112.725 164.035 112.985 164.295 ;
        RECT 112.405 161.755 112.665 162.015 ;
        RECT 112.725 161.755 112.985 162.015 ;
        RECT 109.665 159.475 109.925 159.735 ;
        RECT 109.985 159.475 110.245 159.735 ;
        RECT 111.035 159.475 111.295 159.735 ;
        RECT 111.355 159.475 111.615 159.735 ;
        RECT 112.405 159.475 112.665 159.735 ;
        RECT 112.725 159.475 112.985 159.735 ;
        RECT 109.665 157.195 109.925 157.455 ;
        RECT 109.985 157.195 110.245 157.455 ;
        RECT 111.035 157.195 111.295 157.455 ;
        RECT 111.355 157.195 111.615 157.455 ;
        RECT 112.405 157.195 112.665 157.455 ;
        RECT 112.725 157.195 112.985 157.455 ;
        RECT 109.665 154.915 109.925 155.175 ;
        RECT 109.985 154.915 110.245 155.175 ;
        RECT 111.035 154.915 111.295 155.175 ;
        RECT 111.355 154.915 111.615 155.175 ;
        RECT 112.405 154.915 112.665 155.175 ;
        RECT 112.725 154.915 112.985 155.175 ;
        RECT 109.665 152.635 109.925 152.895 ;
        RECT 109.985 152.635 110.245 152.895 ;
        RECT 111.035 152.635 111.295 152.895 ;
        RECT 111.355 152.635 111.615 152.895 ;
        RECT 112.405 152.635 112.665 152.895 ;
        RECT 112.725 152.635 112.985 152.895 ;
        RECT 109.665 150.355 109.925 150.615 ;
        RECT 109.985 150.355 110.245 150.615 ;
        RECT 111.035 150.355 111.295 150.615 ;
        RECT 111.355 150.355 111.615 150.615 ;
        RECT 112.405 150.355 112.665 150.615 ;
        RECT 112.725 150.355 112.985 150.615 ;
        RECT 109.665 148.075 109.925 148.335 ;
        RECT 109.985 148.075 110.245 148.335 ;
        RECT 111.035 148.075 111.295 148.335 ;
        RECT 111.355 148.075 111.615 148.335 ;
        RECT 112.405 148.075 112.665 148.335 ;
        RECT 112.725 148.075 112.985 148.335 ;
        RECT 109.665 145.795 109.925 146.055 ;
        RECT 109.985 145.795 110.245 146.055 ;
        RECT 111.035 145.795 111.295 146.055 ;
        RECT 111.355 145.795 111.615 146.055 ;
        RECT 112.405 145.795 112.665 146.055 ;
        RECT 112.725 145.795 112.985 146.055 ;
        RECT 109.665 143.515 109.925 143.775 ;
        RECT 109.985 143.515 110.245 143.775 ;
        RECT 111.035 143.515 111.295 143.775 ;
        RECT 111.355 143.515 111.615 143.775 ;
        RECT 112.405 143.515 112.665 143.775 ;
        RECT 112.725 143.515 112.985 143.775 ;
        RECT 109.665 141.235 109.925 141.495 ;
        RECT 109.985 141.235 110.245 141.495 ;
        RECT 111.035 141.235 111.295 141.495 ;
        RECT 111.355 141.235 111.615 141.495 ;
        RECT 112.405 141.235 112.665 141.495 ;
        RECT 112.725 141.235 112.985 141.495 ;
        RECT 109.665 138.955 109.925 139.215 ;
        RECT 109.985 138.955 110.245 139.215 ;
        RECT 111.035 138.955 111.295 139.215 ;
        RECT 111.355 138.955 111.615 139.215 ;
        RECT 112.405 138.955 112.665 139.215 ;
        RECT 112.725 138.955 112.985 139.215 ;
        RECT 109.665 136.675 109.925 136.935 ;
        RECT 109.985 136.675 110.245 136.935 ;
        RECT 109.665 134.395 109.925 134.655 ;
        RECT 109.985 134.395 110.245 134.655 ;
        RECT 109.665 132.115 109.925 132.375 ;
        RECT 109.985 132.115 110.245 132.375 ;
        RECT 109.665 129.835 109.925 130.095 ;
        RECT 109.985 129.835 110.245 130.095 ;
        RECT 109.665 127.555 109.925 127.815 ;
        RECT 109.985 127.555 110.245 127.815 ;
        RECT 109.665 125.275 109.925 125.535 ;
        RECT 109.985 125.275 110.245 125.535 ;
        RECT 109.665 122.995 109.925 123.255 ;
        RECT 109.985 122.995 110.245 123.255 ;
        RECT 109.665 120.715 109.925 120.975 ;
        RECT 109.985 120.715 110.245 120.975 ;
        RECT 109.665 118.435 109.925 118.695 ;
        RECT 109.985 118.435 110.245 118.695 ;
        RECT 109.665 116.155 109.925 116.415 ;
        RECT 109.985 116.155 110.245 116.415 ;
        RECT 109.665 113.875 109.925 114.135 ;
        RECT 109.985 113.875 110.245 114.135 ;
        RECT 109.665 111.595 109.925 111.855 ;
        RECT 109.985 111.595 110.245 111.855 ;
        RECT 109.665 109.315 109.925 109.575 ;
        RECT 109.985 109.315 110.245 109.575 ;
        RECT 109.665 107.035 109.925 107.295 ;
        RECT 109.985 107.035 110.245 107.295 ;
        RECT 109.665 104.755 109.925 105.015 ;
        RECT 109.985 104.755 110.245 105.015 ;
        RECT 109.665 102.475 109.925 102.735 ;
        RECT 109.985 102.475 110.245 102.735 ;
        RECT 109.665 100.195 109.925 100.455 ;
        RECT 109.985 100.195 110.245 100.455 ;
        RECT 109.665 97.915 109.925 98.175 ;
        RECT 109.985 97.915 110.245 98.175 ;
        RECT 109.665 95.635 109.925 95.895 ;
        RECT 109.985 95.635 110.245 95.895 ;
        RECT 109.665 93.355 109.925 93.615 ;
        RECT 109.985 93.355 110.245 93.615 ;
        RECT 109.665 91.075 109.925 91.335 ;
        RECT 109.985 91.075 110.245 91.335 ;
        RECT 109.665 88.795 109.925 89.055 ;
        RECT 109.985 88.795 110.245 89.055 ;
        RECT 109.665 86.515 109.925 86.775 ;
        RECT 109.985 86.515 110.245 86.775 ;
        RECT 109.665 84.235 109.925 84.495 ;
        RECT 109.985 84.235 110.245 84.495 ;
        RECT 109.665 81.955 109.925 82.215 ;
        RECT 109.985 81.955 110.245 82.215 ;
        RECT 109.665 79.675 109.925 79.935 ;
        RECT 109.985 79.675 110.245 79.935 ;
        RECT 109.665 77.395 109.925 77.655 ;
        RECT 109.985 77.395 110.245 77.655 ;
        RECT 109.665 75.115 109.925 75.375 ;
        RECT 109.985 75.115 110.245 75.375 ;
        RECT 109.665 72.835 109.925 73.095 ;
        RECT 109.985 72.835 110.245 73.095 ;
        RECT 109.665 70.555 109.925 70.815 ;
        RECT 109.985 70.555 110.245 70.815 ;
        RECT 111.035 136.675 111.295 136.935 ;
        RECT 111.355 136.675 111.615 136.935 ;
        RECT 111.035 134.395 111.295 134.655 ;
        RECT 111.355 134.395 111.615 134.655 ;
        RECT 111.035 132.115 111.295 132.375 ;
        RECT 111.355 132.115 111.615 132.375 ;
        RECT 111.035 129.835 111.295 130.095 ;
        RECT 111.355 129.835 111.615 130.095 ;
        RECT 111.035 127.555 111.295 127.815 ;
        RECT 111.355 127.555 111.615 127.815 ;
        RECT 111.035 125.275 111.295 125.535 ;
        RECT 111.355 125.275 111.615 125.535 ;
        RECT 111.035 122.995 111.295 123.255 ;
        RECT 111.355 122.995 111.615 123.255 ;
        RECT 111.035 120.715 111.295 120.975 ;
        RECT 111.355 120.715 111.615 120.975 ;
        RECT 111.035 118.435 111.295 118.695 ;
        RECT 111.355 118.435 111.615 118.695 ;
        RECT 111.035 116.155 111.295 116.415 ;
        RECT 111.355 116.155 111.615 116.415 ;
        RECT 111.035 113.875 111.295 114.135 ;
        RECT 111.355 113.875 111.615 114.135 ;
        RECT 111.035 111.595 111.295 111.855 ;
        RECT 111.355 111.595 111.615 111.855 ;
        RECT 111.035 109.315 111.295 109.575 ;
        RECT 111.355 109.315 111.615 109.575 ;
        RECT 111.035 107.035 111.295 107.295 ;
        RECT 111.355 107.035 111.615 107.295 ;
        RECT 111.035 104.755 111.295 105.015 ;
        RECT 111.355 104.755 111.615 105.015 ;
        RECT 111.035 102.475 111.295 102.735 ;
        RECT 111.355 102.475 111.615 102.735 ;
        RECT 111.035 100.195 111.295 100.455 ;
        RECT 111.355 100.195 111.615 100.455 ;
        RECT 112.405 136.675 112.665 136.935 ;
        RECT 112.725 136.675 112.985 136.935 ;
        RECT 112.405 134.395 112.665 134.655 ;
        RECT 112.725 134.395 112.985 134.655 ;
        RECT 112.405 132.115 112.665 132.375 ;
        RECT 112.725 132.115 112.985 132.375 ;
        RECT 112.405 129.835 112.665 130.095 ;
        RECT 112.725 129.835 112.985 130.095 ;
        RECT 112.405 127.555 112.665 127.815 ;
        RECT 112.725 127.555 112.985 127.815 ;
        RECT 112.405 125.275 112.665 125.535 ;
        RECT 112.725 125.275 112.985 125.535 ;
        RECT 112.405 122.995 112.665 123.255 ;
        RECT 112.725 122.995 112.985 123.255 ;
        RECT 112.405 120.715 112.665 120.975 ;
        RECT 112.725 120.715 112.985 120.975 ;
        RECT 112.405 118.435 112.665 118.695 ;
        RECT 112.725 118.435 112.985 118.695 ;
        RECT 112.405 116.155 112.665 116.415 ;
        RECT 112.725 116.155 112.985 116.415 ;
        RECT 112.405 113.875 112.665 114.135 ;
        RECT 112.725 113.875 112.985 114.135 ;
        RECT 122.870 164.665 123.130 164.925 ;
        RECT 123.190 164.665 123.450 164.925 ;
        RECT 124.240 164.665 124.500 164.925 ;
        RECT 124.560 164.665 124.820 164.925 ;
        RECT 115.410 117.075 115.670 117.335 ;
        RECT 115.410 116.755 115.670 117.015 ;
        RECT 115.955 116.620 116.215 116.880 ;
        RECT 116.275 116.620 116.535 116.880 ;
        RECT 115.955 116.190 116.215 116.450 ;
        RECT 116.275 116.190 116.535 116.450 ;
        RECT 115.955 115.760 116.215 116.020 ;
        RECT 116.275 115.760 116.535 116.020 ;
        RECT 122.870 164.035 123.130 164.295 ;
        RECT 123.190 164.035 123.450 164.295 ;
        RECT 123.715 163.885 123.975 164.145 ;
        RECT 124.240 164.035 124.500 164.295 ;
        RECT 124.560 164.035 124.820 164.295 ;
        RECT 123.715 163.565 123.975 163.825 ;
        RECT 123.715 163.245 123.975 163.505 ;
        RECT 123.715 162.925 123.975 163.185 ;
        RECT 123.715 162.605 123.975 162.865 ;
        RECT 123.715 162.285 123.975 162.545 ;
        RECT 122.870 161.755 123.130 162.015 ;
        RECT 123.190 161.755 123.450 162.015 ;
        RECT 123.715 161.965 123.975 162.225 ;
        RECT 123.715 161.645 123.975 161.905 ;
        RECT 124.240 161.755 124.500 162.015 ;
        RECT 124.560 161.755 124.820 162.015 ;
        RECT 123.715 161.325 123.975 161.585 ;
        RECT 123.715 161.005 123.975 161.265 ;
        RECT 123.715 160.685 123.975 160.945 ;
        RECT 123.715 160.365 123.975 160.625 ;
        RECT 123.715 160.045 123.975 160.305 ;
        RECT 122.870 159.475 123.130 159.735 ;
        RECT 123.190 159.475 123.450 159.735 ;
        RECT 123.715 159.725 123.975 159.985 ;
        RECT 123.715 159.405 123.975 159.665 ;
        RECT 124.240 159.475 124.500 159.735 ;
        RECT 124.560 159.475 124.820 159.735 ;
        RECT 123.715 159.085 123.975 159.345 ;
        RECT 123.715 158.765 123.975 159.025 ;
        RECT 123.715 158.445 123.975 158.705 ;
        RECT 123.715 158.125 123.975 158.385 ;
        RECT 123.715 157.805 123.975 158.065 ;
        RECT 123.715 157.485 123.975 157.745 ;
        RECT 122.870 157.195 123.130 157.455 ;
        RECT 123.190 157.195 123.450 157.455 ;
        RECT 123.715 157.165 123.975 157.425 ;
        RECT 124.240 157.195 124.500 157.455 ;
        RECT 124.560 157.195 124.820 157.455 ;
        RECT 123.715 156.845 123.975 157.105 ;
        RECT 123.715 156.525 123.975 156.785 ;
        RECT 123.715 156.205 123.975 156.465 ;
        RECT 123.715 155.885 123.975 156.145 ;
        RECT 123.715 155.565 123.975 155.825 ;
        RECT 123.715 155.245 123.975 155.505 ;
        RECT 122.870 154.915 123.130 155.175 ;
        RECT 123.190 154.915 123.450 155.175 ;
        RECT 123.715 154.925 123.975 155.185 ;
        RECT 124.240 154.915 124.500 155.175 ;
        RECT 124.560 154.915 124.820 155.175 ;
        RECT 123.715 154.605 123.975 154.865 ;
        RECT 123.715 154.285 123.975 154.545 ;
        RECT 123.715 153.965 123.975 154.225 ;
        RECT 123.715 153.645 123.975 153.905 ;
        RECT 123.715 153.325 123.975 153.585 ;
        RECT 123.715 153.005 123.975 153.265 ;
        RECT 122.870 152.635 123.130 152.895 ;
        RECT 123.190 152.635 123.450 152.895 ;
        RECT 123.715 152.685 123.975 152.945 ;
        RECT 124.240 152.635 124.500 152.895 ;
        RECT 124.560 152.635 124.820 152.895 ;
        RECT 123.715 152.365 123.975 152.625 ;
        RECT 123.715 152.045 123.975 152.305 ;
        RECT 123.715 151.725 123.975 151.985 ;
        RECT 123.715 151.405 123.975 151.665 ;
        RECT 123.715 151.085 123.975 151.345 ;
        RECT 123.715 150.765 123.975 151.025 ;
        RECT 122.870 150.355 123.130 150.615 ;
        RECT 123.190 150.355 123.450 150.615 ;
        RECT 123.715 150.445 123.975 150.705 ;
        RECT 123.715 150.125 123.975 150.385 ;
        RECT 124.240 150.355 124.500 150.615 ;
        RECT 124.560 150.355 124.820 150.615 ;
        RECT 123.715 149.805 123.975 150.065 ;
        RECT 123.715 149.485 123.975 149.745 ;
        RECT 123.715 149.165 123.975 149.425 ;
        RECT 123.715 148.845 123.975 149.105 ;
        RECT 123.715 148.525 123.975 148.785 ;
        RECT 122.870 148.075 123.130 148.335 ;
        RECT 123.190 148.075 123.450 148.335 ;
        RECT 123.715 148.205 123.975 148.465 ;
        RECT 123.715 147.885 123.975 148.145 ;
        RECT 124.240 148.075 124.500 148.335 ;
        RECT 124.560 148.075 124.820 148.335 ;
        RECT 123.715 147.565 123.975 147.825 ;
        RECT 123.715 147.245 123.975 147.505 ;
        RECT 123.715 146.925 123.975 147.185 ;
        RECT 123.715 146.605 123.975 146.865 ;
        RECT 123.715 146.285 123.975 146.545 ;
        RECT 122.870 145.795 123.130 146.055 ;
        RECT 123.190 145.795 123.450 146.055 ;
        RECT 123.715 145.965 123.975 146.225 ;
        RECT 123.715 145.645 123.975 145.905 ;
        RECT 124.240 145.795 124.500 146.055 ;
        RECT 124.560 145.795 124.820 146.055 ;
        RECT 123.715 145.325 123.975 145.585 ;
        RECT 123.715 145.005 123.975 145.265 ;
        RECT 123.715 144.685 123.975 144.945 ;
        RECT 123.715 144.365 123.975 144.625 ;
        RECT 123.715 144.045 123.975 144.305 ;
        RECT 122.870 143.515 123.130 143.775 ;
        RECT 123.190 143.515 123.450 143.775 ;
        RECT 123.715 143.725 123.975 143.985 ;
        RECT 123.715 143.405 123.975 143.665 ;
        RECT 124.240 143.515 124.500 143.775 ;
        RECT 124.560 143.515 124.820 143.775 ;
        RECT 123.715 143.085 123.975 143.345 ;
        RECT 123.715 142.765 123.975 143.025 ;
        RECT 123.715 142.445 123.975 142.705 ;
        RECT 123.715 142.125 123.975 142.385 ;
        RECT 123.715 141.805 123.975 142.065 ;
        RECT 122.870 141.235 123.130 141.495 ;
        RECT 123.190 141.235 123.450 141.495 ;
        RECT 123.715 141.485 123.975 141.745 ;
        RECT 123.715 141.165 123.975 141.425 ;
        RECT 124.240 141.235 124.500 141.495 ;
        RECT 124.560 141.235 124.820 141.495 ;
        RECT 123.715 140.845 123.975 141.105 ;
        RECT 123.715 140.525 123.975 140.785 ;
        RECT 123.715 140.205 123.975 140.465 ;
        RECT 123.715 139.885 123.975 140.145 ;
        RECT 123.715 139.565 123.975 139.825 ;
        RECT 123.715 139.245 123.975 139.505 ;
        RECT 122.870 138.955 123.130 139.215 ;
        RECT 123.190 138.955 123.450 139.215 ;
        RECT 123.715 138.925 123.975 139.185 ;
        RECT 124.240 138.955 124.500 139.215 ;
        RECT 124.560 138.955 124.820 139.215 ;
        RECT 123.715 138.605 123.975 138.865 ;
        RECT 123.715 138.285 123.975 138.545 ;
        RECT 123.715 137.965 123.975 138.225 ;
        RECT 123.715 137.645 123.975 137.905 ;
        RECT 123.715 137.325 123.975 137.585 ;
        RECT 123.715 137.005 123.975 137.265 ;
        RECT 122.870 136.675 123.130 136.935 ;
        RECT 123.190 136.675 123.450 136.935 ;
        RECT 123.715 136.685 123.975 136.945 ;
        RECT 122.870 134.395 123.130 134.655 ;
        RECT 123.190 134.395 123.450 134.655 ;
        RECT 122.870 132.115 123.130 132.375 ;
        RECT 123.190 132.115 123.450 132.375 ;
        RECT 122.870 129.835 123.130 130.095 ;
        RECT 123.190 129.835 123.450 130.095 ;
        RECT 122.870 127.555 123.130 127.815 ;
        RECT 123.190 127.555 123.450 127.815 ;
        RECT 122.870 125.275 123.130 125.535 ;
        RECT 123.190 125.275 123.450 125.535 ;
        RECT 122.870 122.995 123.130 123.255 ;
        RECT 123.190 122.995 123.450 123.255 ;
        RECT 122.870 120.715 123.130 120.975 ;
        RECT 123.190 120.715 123.450 120.975 ;
        RECT 122.870 118.435 123.130 118.695 ;
        RECT 123.190 118.435 123.450 118.695 ;
        RECT 122.870 116.155 123.130 116.415 ;
        RECT 123.190 116.155 123.450 116.415 ;
        RECT 119.215 114.235 119.475 114.495 ;
        RECT 119.535 114.235 119.795 114.495 ;
        RECT 119.855 114.235 120.115 114.495 ;
        RECT 120.390 114.130 120.650 114.390 ;
        RECT 112.405 111.595 112.665 111.855 ;
        RECT 112.725 111.595 112.985 111.855 ;
        RECT 115.955 111.950 116.215 112.210 ;
        RECT 116.275 111.950 116.535 112.210 ;
        RECT 112.405 109.315 112.665 109.575 ;
        RECT 112.725 109.315 112.985 109.575 ;
        RECT 112.405 107.035 112.665 107.295 ;
        RECT 112.725 107.035 112.985 107.295 ;
        RECT 112.405 104.755 112.665 105.015 ;
        RECT 112.725 104.755 112.985 105.015 ;
        RECT 112.405 102.475 112.665 102.735 ;
        RECT 112.725 102.475 112.985 102.735 ;
        RECT 112.405 100.195 112.665 100.455 ;
        RECT 112.725 100.195 112.985 100.455 ;
        RECT 111.880 99.495 112.140 99.755 ;
        RECT 111.880 99.175 112.140 99.435 ;
        RECT 111.880 98.855 112.140 99.115 ;
        RECT 111.880 98.535 112.140 98.795 ;
        RECT 111.035 97.915 111.295 98.175 ;
        RECT 111.355 97.915 111.615 98.175 ;
        RECT 111.035 95.635 111.295 95.895 ;
        RECT 111.355 95.635 111.615 95.895 ;
        RECT 111.035 93.355 111.295 93.615 ;
        RECT 111.355 93.355 111.615 93.615 ;
        RECT 111.035 91.075 111.295 91.335 ;
        RECT 111.355 91.075 111.615 91.335 ;
        RECT 111.035 88.795 111.295 89.055 ;
        RECT 111.355 88.795 111.615 89.055 ;
        RECT 111.035 86.515 111.295 86.775 ;
        RECT 111.355 86.515 111.615 86.775 ;
        RECT 111.035 84.235 111.295 84.495 ;
        RECT 111.355 84.235 111.615 84.495 ;
        RECT 111.035 81.955 111.295 82.215 ;
        RECT 111.355 81.955 111.615 82.215 ;
        RECT 111.035 79.675 111.295 79.935 ;
        RECT 111.355 79.675 111.615 79.935 ;
        RECT 111.035 77.395 111.295 77.655 ;
        RECT 111.355 77.395 111.615 77.655 ;
        RECT 111.035 75.115 111.295 75.375 ;
        RECT 111.355 75.115 111.615 75.375 ;
        RECT 111.035 72.835 111.295 73.095 ;
        RECT 111.355 72.835 111.615 73.095 ;
        RECT 111.035 70.555 111.295 70.815 ;
        RECT 111.355 70.555 111.615 70.815 ;
        RECT 112.405 97.915 112.665 98.175 ;
        RECT 112.725 97.915 112.985 98.175 ;
        RECT 112.405 95.635 112.665 95.895 ;
        RECT 112.725 95.635 112.985 95.895 ;
        RECT 112.405 93.355 112.665 93.615 ;
        RECT 112.725 93.355 112.985 93.615 ;
        RECT 112.405 91.075 112.665 91.335 ;
        RECT 112.725 91.075 112.985 91.335 ;
        RECT 112.405 88.795 112.665 89.055 ;
        RECT 112.725 88.795 112.985 89.055 ;
        RECT 112.405 86.515 112.665 86.775 ;
        RECT 112.725 86.515 112.985 86.775 ;
        RECT 112.405 84.235 112.665 84.495 ;
        RECT 112.725 84.235 112.985 84.495 ;
        RECT 112.405 81.955 112.665 82.215 ;
        RECT 112.725 81.955 112.985 82.215 ;
        RECT 112.405 79.675 112.665 79.935 ;
        RECT 112.725 79.675 112.985 79.935 ;
        RECT 115.955 111.520 116.215 111.780 ;
        RECT 116.275 111.520 116.535 111.780 ;
        RECT 115.955 111.090 116.215 111.350 ;
        RECT 116.275 111.090 116.535 111.350 ;
        RECT 116.820 110.525 117.080 110.785 ;
        RECT 116.820 110.205 117.080 110.465 ;
        RECT 120.390 113.810 120.650 114.070 ;
        RECT 119.215 113.375 119.475 113.635 ;
        RECT 119.535 113.375 119.795 113.635 ;
        RECT 119.855 113.375 120.115 113.635 ;
        RECT 120.390 113.490 120.650 113.750 ;
        RECT 122.870 113.875 123.130 114.135 ;
        RECT 123.190 113.875 123.450 114.135 ;
        RECT 115.410 82.875 115.670 83.135 ;
        RECT 115.410 82.555 115.670 82.815 ;
        RECT 115.955 82.420 116.215 82.680 ;
        RECT 116.275 82.420 116.535 82.680 ;
        RECT 115.955 81.990 116.215 82.250 ;
        RECT 116.275 81.990 116.535 82.250 ;
        RECT 115.955 81.560 116.215 81.820 ;
        RECT 116.275 81.560 116.535 81.820 ;
        RECT 119.215 80.035 119.475 80.295 ;
        RECT 119.535 80.035 119.795 80.295 ;
        RECT 119.855 80.035 120.115 80.295 ;
        RECT 120.390 79.930 120.650 80.190 ;
        RECT 112.405 77.395 112.665 77.655 ;
        RECT 112.725 77.395 112.985 77.655 ;
        RECT 115.955 77.750 116.215 78.010 ;
        RECT 116.275 77.750 116.535 78.010 ;
        RECT 112.405 75.115 112.665 75.375 ;
        RECT 112.725 75.115 112.985 75.375 ;
        RECT 112.405 72.835 112.665 73.095 ;
        RECT 112.725 72.835 112.985 73.095 ;
        RECT 112.405 70.555 112.665 70.815 ;
        RECT 112.725 70.555 112.985 70.815 ;
        RECT 111.880 69.740 112.140 70.000 ;
        RECT 111.880 69.420 112.140 69.680 ;
        RECT 111.880 69.100 112.140 69.360 ;
        RECT 109.665 68.275 109.925 68.535 ;
        RECT 109.985 68.275 110.245 68.535 ;
        RECT 111.035 68.275 111.295 68.535 ;
        RECT 111.355 68.275 111.615 68.535 ;
        RECT 112.405 68.275 112.665 68.535 ;
        RECT 112.725 68.275 112.985 68.535 ;
        RECT 109.665 65.995 109.925 66.255 ;
        RECT 109.985 65.995 110.245 66.255 ;
        RECT 109.665 63.715 109.925 63.975 ;
        RECT 109.985 63.715 110.245 63.975 ;
        RECT 111.035 65.995 111.295 66.255 ;
        RECT 111.355 65.995 111.615 66.255 ;
        RECT 111.035 63.715 111.295 63.975 ;
        RECT 111.355 63.715 111.615 63.975 ;
        RECT 112.405 65.995 112.665 66.255 ;
        RECT 112.725 65.995 112.985 66.255 ;
        RECT 112.405 63.715 112.665 63.975 ;
        RECT 112.725 63.715 112.985 63.975 ;
        RECT 115.955 77.320 116.215 77.580 ;
        RECT 116.275 77.320 116.535 77.580 ;
        RECT 115.955 76.890 116.215 77.150 ;
        RECT 116.275 76.890 116.535 77.150 ;
        RECT 116.820 76.325 117.080 76.585 ;
        RECT 116.820 76.005 117.080 76.265 ;
        RECT 115.805 75.360 116.065 75.620 ;
        RECT 116.125 75.360 116.385 75.620 ;
        RECT 120.390 79.610 120.650 79.870 ;
        RECT 119.215 79.175 119.475 79.435 ;
        RECT 119.535 79.175 119.795 79.435 ;
        RECT 119.855 79.175 120.115 79.435 ;
        RECT 120.390 79.290 120.650 79.550 ;
        RECT 122.870 111.595 123.130 111.855 ;
        RECT 123.190 111.595 123.450 111.855 ;
        RECT 122.870 109.315 123.130 109.575 ;
        RECT 123.190 109.315 123.450 109.575 ;
        RECT 122.870 107.035 123.130 107.295 ;
        RECT 123.190 107.035 123.450 107.295 ;
        RECT 122.870 104.755 123.130 105.015 ;
        RECT 123.190 104.755 123.450 105.015 ;
        RECT 122.870 102.475 123.130 102.735 ;
        RECT 123.190 102.475 123.450 102.735 ;
        RECT 122.870 100.195 123.130 100.455 ;
        RECT 123.190 100.195 123.450 100.455 ;
        RECT 122.870 97.915 123.130 98.175 ;
        RECT 123.190 97.915 123.450 98.175 ;
        RECT 122.870 95.635 123.130 95.895 ;
        RECT 123.190 95.635 123.450 95.895 ;
        RECT 122.870 93.355 123.130 93.615 ;
        RECT 123.190 93.355 123.450 93.615 ;
        RECT 122.870 91.075 123.130 91.335 ;
        RECT 123.190 91.075 123.450 91.335 ;
        RECT 122.870 88.795 123.130 89.055 ;
        RECT 123.190 88.795 123.450 89.055 ;
        RECT 122.870 86.515 123.130 86.775 ;
        RECT 123.190 86.515 123.450 86.775 ;
        RECT 122.870 84.235 123.130 84.495 ;
        RECT 123.190 84.235 123.450 84.495 ;
        RECT 122.345 83.410 122.605 83.670 ;
        RECT 122.345 83.090 122.605 83.350 ;
        RECT 122.345 82.770 122.605 83.030 ;
        RECT 124.240 136.675 124.500 136.935 ;
        RECT 124.560 136.675 124.820 136.935 ;
        RECT 124.240 134.395 124.500 134.655 ;
        RECT 124.560 134.395 124.820 134.655 ;
        RECT 124.240 132.115 124.500 132.375 ;
        RECT 124.560 132.115 124.820 132.375 ;
        RECT 124.240 129.835 124.500 130.095 ;
        RECT 124.560 129.835 124.820 130.095 ;
        RECT 124.240 127.555 124.500 127.815 ;
        RECT 124.560 127.555 124.820 127.815 ;
        RECT 124.240 125.275 124.500 125.535 ;
        RECT 124.560 125.275 124.820 125.535 ;
        RECT 124.240 122.995 124.500 123.255 ;
        RECT 124.560 122.995 124.820 123.255 ;
        RECT 124.240 120.715 124.500 120.975 ;
        RECT 124.560 120.715 124.820 120.975 ;
        RECT 124.240 118.435 124.500 118.695 ;
        RECT 124.560 118.435 124.820 118.695 ;
        RECT 124.240 116.155 124.500 116.415 ;
        RECT 124.560 116.155 124.820 116.415 ;
        RECT 124.240 113.875 124.500 114.135 ;
        RECT 124.560 113.875 124.820 114.135 ;
        RECT 124.240 111.595 124.500 111.855 ;
        RECT 124.560 111.595 124.820 111.855 ;
        RECT 124.240 109.315 124.500 109.575 ;
        RECT 124.560 109.315 124.820 109.575 ;
        RECT 124.240 107.035 124.500 107.295 ;
        RECT 124.560 107.035 124.820 107.295 ;
        RECT 124.240 104.755 124.500 105.015 ;
        RECT 124.560 104.755 124.820 105.015 ;
        RECT 124.240 102.475 124.500 102.735 ;
        RECT 124.560 102.475 124.820 102.735 ;
        RECT 124.240 100.195 124.500 100.455 ;
        RECT 124.560 100.195 124.820 100.455 ;
        RECT 124.240 97.915 124.500 98.175 ;
        RECT 124.560 97.915 124.820 98.175 ;
        RECT 124.240 95.635 124.500 95.895 ;
        RECT 124.560 95.635 124.820 95.895 ;
        RECT 124.240 93.355 124.500 93.615 ;
        RECT 124.560 93.355 124.820 93.615 ;
        RECT 124.240 91.075 124.500 91.335 ;
        RECT 124.560 91.075 124.820 91.335 ;
        RECT 124.240 88.795 124.500 89.055 ;
        RECT 124.560 88.795 124.820 89.055 ;
        RECT 124.240 86.515 124.500 86.775 ;
        RECT 124.560 86.515 124.820 86.775 ;
        RECT 124.240 84.235 124.500 84.495 ;
        RECT 124.560 84.235 124.820 84.495 ;
        RECT 123.715 83.410 123.975 83.670 ;
        RECT 123.715 83.090 123.975 83.350 ;
        RECT 123.715 82.770 123.975 83.030 ;
        RECT 122.870 81.955 123.130 82.215 ;
        RECT 123.190 81.955 123.450 82.215 ;
        RECT 124.240 81.955 124.500 82.215 ;
        RECT 124.560 81.955 124.820 82.215 ;
        RECT 122.870 79.675 123.130 79.935 ;
        RECT 123.190 79.675 123.450 79.935 ;
        RECT 124.240 79.675 124.500 79.935 ;
        RECT 124.560 79.675 124.820 79.935 ;
        RECT 122.870 77.395 123.130 77.655 ;
        RECT 123.190 77.395 123.450 77.655 ;
        RECT 124.240 77.395 124.500 77.655 ;
        RECT 124.560 77.395 124.820 77.655 ;
        RECT 122.870 76.765 123.130 77.025 ;
        RECT 123.190 76.765 123.450 77.025 ;
        RECT 124.240 76.765 124.500 77.025 ;
        RECT 124.560 76.765 124.820 77.025 ;
        RECT 109.665 63.045 109.925 63.305 ;
        RECT 109.985 63.045 110.245 63.305 ;
        RECT 111.035 63.045 111.295 63.305 ;
        RECT 111.355 63.045 111.615 63.305 ;
        RECT 112.405 63.045 112.665 63.305 ;
        RECT 112.725 63.045 112.985 63.305 ;
        RECT 115.805 70.585 116.065 70.845 ;
        RECT 116.125 70.585 116.385 70.845 ;
        RECT 115.805 69.915 116.065 70.175 ;
        RECT 116.125 69.915 116.385 70.175 ;
        RECT 115.260 69.430 115.520 69.690 ;
        RECT 115.260 69.110 115.520 69.370 ;
        RECT 115.260 68.790 115.520 69.050 ;
        RECT 119.500 70.305 119.760 70.565 ;
        RECT 119.820 70.305 120.080 70.565 ;
        RECT 119.500 69.635 119.760 69.895 ;
        RECT 119.820 69.635 120.080 69.895 ;
        RECT 120.365 69.720 120.625 69.980 ;
        RECT 119.500 69.205 119.760 69.465 ;
        RECT 119.820 69.205 120.080 69.465 ;
        RECT 120.365 69.400 120.625 69.660 ;
        RECT 119.500 68.775 119.760 69.035 ;
        RECT 119.820 68.775 120.080 69.035 ;
        RECT 119.500 68.360 119.760 68.620 ;
        RECT 119.820 68.360 120.080 68.620 ;
        RECT 115.805 67.635 116.065 67.895 ;
        RECT 116.125 67.635 116.385 67.895 ;
        RECT 115.805 65.355 116.065 65.615 ;
        RECT 116.125 65.355 116.385 65.615 ;
        RECT 115.805 63.075 116.065 63.335 ;
        RECT 116.125 63.075 116.385 63.335 ;
        RECT 115.805 60.795 116.065 61.055 ;
        RECT 116.125 60.795 116.385 61.055 ;
        RECT 119.500 67.915 119.760 68.175 ;
        RECT 119.820 67.915 120.080 68.175 ;
        RECT 119.500 67.500 119.760 67.760 ;
        RECT 119.820 67.500 120.080 67.760 ;
        RECT 123.080 69.730 123.340 69.990 ;
        RECT 123.080 69.410 123.340 69.670 ;
        RECT 123.080 69.090 123.340 69.350 ;
        RECT 122.215 68.775 122.475 69.035 ;
        RECT 122.535 68.775 122.795 69.035 ;
        RECT 122.215 68.345 122.475 68.605 ;
        RECT 122.535 68.345 122.795 68.605 ;
        RECT 122.215 67.915 122.475 68.175 ;
        RECT 122.535 67.915 122.795 68.175 ;
        RECT 122.215 67.485 122.475 67.745 ;
        RECT 122.535 67.485 122.795 67.745 ;
        RECT 119.500 67.055 119.760 67.315 ;
        RECT 119.820 67.055 120.080 67.315 ;
        RECT 122.215 67.055 122.475 67.315 ;
        RECT 122.535 67.055 122.795 67.315 ;
        RECT 119.500 66.625 119.760 66.885 ;
        RECT 119.820 66.625 120.080 66.885 ;
        RECT 119.500 66.195 119.760 66.455 ;
        RECT 119.820 66.195 120.080 66.455 ;
        RECT 125.485 70.265 125.745 70.525 ;
        RECT 125.805 70.265 126.065 70.525 ;
        RECT 115.805 60.125 116.065 60.385 ;
        RECT 116.125 60.125 116.385 60.385 ;
        RECT 119.500 64.385 119.760 64.645 ;
        RECT 119.820 64.385 120.080 64.645 ;
        RECT 120.475 64.360 120.735 64.620 ;
        RECT 119.500 63.955 119.760 64.215 ;
        RECT 119.820 63.955 120.080 64.215 ;
        RECT 120.475 64.040 120.735 64.300 ;
        RECT 119.500 63.525 119.760 63.785 ;
        RECT 119.820 63.525 120.080 63.785 ;
        RECT 120.475 63.720 120.735 63.980 ;
        RECT 119.500 63.110 119.760 63.370 ;
        RECT 119.820 63.110 120.080 63.370 ;
        RECT 119.500 62.665 119.760 62.925 ;
        RECT 119.820 62.665 120.080 62.925 ;
        RECT 119.500 62.250 119.760 62.510 ;
        RECT 119.820 62.250 120.080 62.510 ;
        RECT 122.215 63.525 122.475 63.785 ;
        RECT 122.535 63.525 122.795 63.785 ;
        RECT 125.485 69.635 125.745 69.895 ;
        RECT 125.805 69.635 126.065 69.895 ;
        RECT 125.485 69.205 125.745 69.465 ;
        RECT 125.805 69.205 126.065 69.465 ;
        RECT 125.485 68.775 125.745 69.035 ;
        RECT 125.805 68.775 126.065 69.035 ;
        RECT 125.485 68.345 125.745 68.605 ;
        RECT 125.805 68.345 126.065 68.605 ;
        RECT 125.485 67.915 125.745 68.175 ;
        RECT 125.805 67.915 126.065 68.175 ;
        RECT 125.485 67.485 125.745 67.745 ;
        RECT 125.805 67.485 126.065 67.745 ;
        RECT 125.485 67.055 125.745 67.315 ;
        RECT 125.805 67.055 126.065 67.315 ;
        RECT 125.485 66.625 125.745 66.885 ;
        RECT 125.805 66.625 126.065 66.885 ;
        RECT 125.485 66.195 125.745 66.455 ;
        RECT 125.805 66.195 126.065 66.455 ;
        RECT 125.485 65.765 125.745 66.025 ;
        RECT 125.805 65.765 126.065 66.025 ;
        RECT 126.335 65.640 126.595 65.900 ;
        RECT 125.485 65.335 125.745 65.595 ;
        RECT 125.805 65.335 126.065 65.595 ;
        RECT 126.335 65.320 126.595 65.580 ;
        RECT 125.485 64.905 125.745 65.165 ;
        RECT 125.805 64.905 126.065 65.165 ;
        RECT 126.335 65.000 126.595 65.260 ;
        RECT 125.485 64.475 125.745 64.735 ;
        RECT 125.805 64.475 126.065 64.735 ;
        RECT 122.215 63.095 122.475 63.355 ;
        RECT 122.535 63.095 122.795 63.355 ;
        RECT 122.215 62.665 122.475 62.925 ;
        RECT 122.535 62.665 122.795 62.925 ;
        RECT 122.215 62.235 122.475 62.495 ;
        RECT 122.535 62.235 122.795 62.495 ;
        RECT 119.500 61.805 119.760 62.065 ;
        RECT 119.820 61.805 120.080 62.065 ;
        RECT 122.215 61.805 122.475 62.065 ;
        RECT 122.535 61.805 122.795 62.065 ;
        RECT 119.500 61.375 119.760 61.635 ;
        RECT 119.820 61.375 120.080 61.635 ;
        RECT 119.500 60.945 119.760 61.205 ;
        RECT 119.820 60.945 120.080 61.205 ;
        RECT 123.080 61.420 123.340 61.680 ;
        RECT 123.080 61.100 123.340 61.360 ;
        RECT 119.500 60.315 119.760 60.575 ;
        RECT 119.820 60.315 120.080 60.575 ;
        RECT 125.485 64.045 125.745 64.305 ;
        RECT 125.805 64.045 126.065 64.305 ;
        RECT 125.485 63.615 125.745 63.875 ;
        RECT 125.805 63.615 126.065 63.875 ;
        RECT 125.485 63.185 125.745 63.445 ;
        RECT 125.805 63.185 126.065 63.445 ;
        RECT 125.485 62.755 125.745 63.015 ;
        RECT 125.805 62.755 126.065 63.015 ;
        RECT 125.485 62.325 125.745 62.585 ;
        RECT 125.805 62.325 126.065 62.585 ;
        RECT 125.485 61.895 125.745 62.155 ;
        RECT 125.805 61.895 126.065 62.155 ;
        RECT 125.485 61.465 125.745 61.725 ;
        RECT 125.805 61.465 126.065 61.725 ;
        RECT 125.485 61.035 125.745 61.295 ;
        RECT 125.805 61.035 126.065 61.295 ;
        RECT 125.485 60.405 125.745 60.665 ;
        RECT 125.805 60.405 126.065 60.665 ;
      LAYER met2 ;
        RECT 127.375 211.800 144.155 212.130 ;
        RECT 115.355 210.970 158.265 211.300 ;
        RECT 120.335 210.140 147.830 210.470 ;
        RECT 157.665 210.220 158.265 210.970 ;
        RECT 123.680 209.040 157.165 209.640 ;
        RECT 156.565 208.960 157.165 209.040 ;
        RECT 117.715 207.940 142.530 208.540 ;
        RECT 106.100 206.445 118.065 207.045 ;
        RECT 117.695 205.965 118.065 206.445 ;
        RECT 84.950 174.320 85.250 174.890 ;
        RECT 45.995 173.720 85.250 174.320 ;
        RECT 108.195 173.840 109.195 174.130 ;
        RECT 112.045 173.840 113.045 174.130 ;
        RECT 45.995 15.375 46.595 173.720 ;
        RECT 88.630 173.220 88.930 173.790 ;
        RECT 47.095 172.620 88.930 173.220 ;
        RECT 108.195 173.175 109.195 173.455 ;
        RECT 108.195 172.745 109.195 173.025 ;
        RECT 110.205 172.675 110.535 173.445 ;
        RECT 112.045 173.175 113.045 173.455 ;
        RECT 112.045 172.745 113.045 173.025 ;
        RECT 47.095 16.475 47.695 172.620 ;
        RECT 108.195 172.315 109.195 172.595 ;
        RECT 112.045 172.315 113.045 172.595 ;
        RECT 108.195 171.885 113.545 172.165 ;
        RECT 108.195 171.455 109.195 171.735 ;
        RECT 110.205 171.305 110.535 171.885 ;
        RECT 112.045 171.455 113.045 171.735 ;
        RECT 108.195 171.025 113.545 171.305 ;
        RECT 108.195 170.595 109.195 170.875 ;
        RECT 110.205 170.670 110.535 171.025 ;
        RECT 108.195 170.165 109.195 170.445 ;
        RECT 108.195 169.735 109.195 170.015 ;
        RECT 110.195 169.790 110.535 170.670 ;
        RECT 112.045 170.595 113.045 170.875 ;
        RECT 112.045 170.165 113.045 170.445 ;
        RECT 108.195 169.060 109.195 169.350 ;
        RECT 110.195 167.605 110.525 169.790 ;
        RECT 112.045 169.735 113.045 170.015 ;
        RECT 112.045 169.060 113.045 169.350 ;
        RECT 116.785 167.605 117.115 168.025 ;
        RECT 110.195 167.275 117.115 167.605 ;
        RECT 116.785 166.855 117.115 167.275 ;
        RECT 109.605 164.690 110.305 164.980 ;
        RECT 110.975 164.690 111.675 164.980 ;
        RECT 112.345 164.690 113.045 164.980 ;
        RECT 122.810 164.650 123.510 164.940 ;
        RECT 109.605 164.025 110.305 164.305 ;
        RECT 110.975 164.025 111.675 164.305 ;
        RECT 112.345 164.025 113.045 164.305 ;
        RECT 122.810 164.025 123.510 164.305 ;
        RECT 109.605 161.745 110.305 162.025 ;
        RECT 110.975 161.745 111.675 162.025 ;
        RECT 112.345 161.745 113.045 162.025 ;
        RECT 122.810 161.745 123.510 162.025 ;
        RECT 123.680 159.745 124.010 166.580 ;
        RECT 124.180 164.650 124.880 164.940 ;
        RECT 124.180 164.025 124.880 164.305 ;
        RECT 124.180 161.745 124.880 162.025 ;
        RECT 109.605 159.465 110.305 159.745 ;
        RECT 110.975 159.465 111.675 159.745 ;
        RECT 112.345 159.465 113.045 159.745 ;
        RECT 122.810 159.465 124.880 159.745 ;
        RECT 109.605 157.185 113.045 157.465 ;
        RECT 122.810 157.185 123.510 157.465 ;
        RECT 109.605 154.905 110.305 155.185 ;
        RECT 78.045 154.200 106.700 154.800 ;
        RECT 78.045 153.100 106.700 153.700 ;
        RECT 106.100 152.620 106.700 153.100 ;
        RECT 110.475 152.905 110.805 157.185 ;
        RECT 110.975 154.905 111.675 155.185 ;
        RECT 111.845 152.905 112.175 157.185 ;
        RECT 123.680 155.185 124.010 159.465 ;
        RECT 124.180 157.185 124.880 157.465 ;
        RECT 112.345 154.905 113.045 155.185 ;
        RECT 122.810 154.905 124.880 155.185 ;
        RECT 109.605 152.625 113.045 152.905 ;
        RECT 122.810 152.625 123.510 152.905 ;
        RECT 63.150 151.930 71.640 152.210 ;
        RECT 57.150 151.440 58.150 151.730 ;
        RECT 60.740 151.440 61.740 151.730 ;
        RECT 65.405 151.440 65.905 151.730 ;
        RECT 60.740 150.775 61.740 151.055 ;
        RECT 65.405 150.775 65.905 151.055 ;
        RECT 71.310 151.040 71.640 151.930 ;
        RECT 87.150 151.930 95.640 152.210 ;
        RECT 87.150 151.040 87.480 151.930 ;
        RECT 92.885 151.440 93.385 151.730 ;
        RECT 97.050 151.440 98.050 151.730 ;
        RECT 100.640 151.440 101.640 151.730 ;
        RECT 92.885 150.775 93.385 151.055 ;
        RECT 97.050 150.775 98.050 151.055 ;
        RECT 109.605 150.345 110.305 150.625 ;
        RECT 60.740 149.995 61.740 150.275 ;
        RECT 65.405 149.995 65.905 150.275 ;
        RECT 92.885 149.995 93.385 150.275 ;
        RECT 97.050 149.995 98.050 150.275 ;
        RECT 60.740 149.215 61.740 149.495 ;
        RECT 63.170 149.050 63.500 149.930 ;
        RECT 65.405 149.215 65.905 149.495 ;
        RECT 92.885 149.215 93.385 149.495 ;
        RECT 61.930 148.760 63.500 149.050 ;
        RECT 95.290 149.050 95.620 149.930 ;
        RECT 97.050 149.215 98.050 149.495 ;
        RECT 95.290 148.760 96.860 149.050 ;
        RECT 61.930 148.150 62.260 148.760 ;
        RECT 96.530 148.150 96.860 148.760 ;
        RECT 110.475 148.345 110.805 152.625 ;
        RECT 110.975 150.345 111.675 150.625 ;
        RECT 111.845 148.345 112.175 152.625 ;
        RECT 123.680 150.625 124.010 154.905 ;
        RECT 124.180 152.625 124.880 152.905 ;
        RECT 112.345 150.345 113.045 150.625 ;
        RECT 122.810 150.345 124.880 150.625 ;
        RECT 109.605 148.065 113.045 148.345 ;
        RECT 122.810 148.065 123.510 148.345 ;
        RECT 64.885 147.215 65.215 147.525 ;
        RECT 93.575 147.215 93.905 147.525 ;
        RECT 60.740 146.935 63.435 147.215 ;
        RECT 63.765 146.935 65.215 147.215 ;
        RECT 65.405 146.935 72.465 147.215 ;
        RECT 63.765 146.045 64.095 146.935 ;
        RECT 64.885 146.625 65.215 146.935 ;
        RECT 72.135 146.045 72.465 146.935 ;
        RECT 86.325 146.935 93.385 147.215 ;
        RECT 93.575 146.935 95.025 147.215 ;
        RECT 95.355 146.935 98.050 147.215 ;
        RECT 86.325 146.045 86.655 146.935 ;
        RECT 93.575 146.625 93.905 146.935 ;
        RECT 94.695 146.045 95.025 146.935 ;
        RECT 109.605 145.785 110.305 146.065 ;
        RECT 60.740 144.655 61.740 144.935 ;
        RECT 65.405 144.655 65.905 144.935 ;
        RECT 92.885 144.655 93.385 144.935 ;
        RECT 97.050 144.655 98.050 144.935 ;
        RECT 60.740 143.875 61.740 144.155 ;
        RECT 65.405 143.875 65.905 144.155 ;
        RECT 92.885 143.875 93.385 144.155 ;
        RECT 97.050 143.875 98.050 144.155 ;
        RECT 110.475 143.785 110.805 148.065 ;
        RECT 110.975 145.785 111.675 146.065 ;
        RECT 111.845 143.785 112.175 148.065 ;
        RECT 123.680 146.065 124.010 150.345 ;
        RECT 124.180 148.065 124.880 148.345 ;
        RECT 112.345 145.785 113.045 146.065 ;
        RECT 122.810 145.785 124.880 146.065 ;
        RECT 109.605 143.505 113.045 143.785 ;
        RECT 122.810 143.505 123.510 143.785 ;
        RECT 60.740 143.095 61.740 143.375 ;
        RECT 65.405 143.095 65.905 143.375 ;
        RECT 92.885 143.095 93.385 143.375 ;
        RECT 97.050 143.095 98.050 143.375 ;
        RECT 73.560 142.720 74.060 143.010 ;
        RECT 76.300 142.720 76.800 143.010 ;
        RECT 81.990 142.720 82.490 143.010 ;
        RECT 84.730 142.720 85.230 143.010 ;
        RECT 60.740 142.315 61.740 142.595 ;
        RECT 65.405 142.420 65.905 142.710 ;
        RECT 92.885 142.420 93.385 142.710 ;
        RECT 73.560 142.095 74.060 142.375 ;
        RECT 57.150 141.535 58.150 141.815 ;
        RECT 59.255 141.535 61.740 141.815 ;
        RECT 76.300 141.695 76.800 141.975 ;
        RECT 57.150 139.255 58.150 139.535 ;
        RECT 59.255 137.255 59.585 141.535 ;
        RECT 78.045 141.370 78.645 142.145 ;
        RECT 61.930 141.040 78.645 141.370 ;
        RECT 80.145 141.370 80.745 142.145 ;
        RECT 84.730 142.095 85.230 142.375 ;
        RECT 97.050 142.315 98.050 142.595 ;
        RECT 81.990 141.695 82.490 141.975 ;
        RECT 97.050 141.535 99.535 141.815 ;
        RECT 100.640 141.535 101.640 141.815 ;
        RECT 80.145 141.040 96.860 141.370 ;
        RECT 61.930 140.470 62.260 141.040 ;
        RECT 73.040 140.790 73.370 141.040 ;
        RECT 85.420 140.790 85.750 141.040 ;
        RECT 96.530 140.470 96.860 141.040 ;
        RECT 75.035 139.815 75.405 140.015 ;
        RECT 73.560 139.535 75.405 139.815 ;
        RECT 60.740 139.255 63.435 139.535 ;
        RECT 75.035 139.335 75.405 139.535 ;
        RECT 83.385 139.815 83.755 140.015 ;
        RECT 83.385 139.535 85.230 139.815 ;
        RECT 83.385 139.335 83.755 139.535 ;
        RECT 95.355 139.255 98.050 139.535 ;
        RECT 65.405 138.230 65.905 138.520 ;
        RECT 69.160 138.230 70.160 138.520 ;
        RECT 76.300 138.415 76.800 138.695 ;
        RECT 81.990 138.415 82.490 138.695 ;
        RECT 88.630 138.230 89.630 138.520 ;
        RECT 92.885 138.230 93.385 138.520 ;
        RECT 65.405 137.565 65.905 137.845 ;
        RECT 69.160 137.565 70.160 137.845 ;
        RECT 88.630 137.565 89.630 137.845 ;
        RECT 92.885 137.565 93.385 137.845 ;
        RECT 72.135 137.255 74.060 137.535 ;
        RECT 84.730 137.255 86.655 137.535 ;
        RECT 99.205 137.255 99.535 141.535 ;
        RECT 109.605 141.225 110.305 141.505 ;
        RECT 100.640 139.255 101.640 139.535 ;
        RECT 110.475 139.225 110.805 143.505 ;
        RECT 110.975 141.225 111.675 141.505 ;
        RECT 111.845 139.225 112.175 143.505 ;
        RECT 123.680 141.505 124.010 145.785 ;
        RECT 124.180 143.505 124.880 143.785 ;
        RECT 112.345 141.225 113.045 141.505 ;
        RECT 122.810 141.225 124.880 141.505 ;
        RECT 109.605 138.945 113.045 139.225 ;
        RECT 122.810 138.945 123.510 139.225 ;
        RECT 57.150 136.975 58.150 137.255 ;
        RECT 59.255 136.975 61.740 137.255 ;
        RECT 57.150 134.695 58.150 134.975 ;
        RECT 59.255 132.695 59.585 136.975 ;
        RECT 65.405 136.285 65.905 136.565 ;
        RECT 69.160 136.285 70.160 136.565 ;
        RECT 65.405 135.005 65.905 135.285 ;
        RECT 69.160 135.005 70.160 135.285 ;
        RECT 60.740 134.695 65.215 134.975 ;
        RECT 64.885 134.075 65.215 134.695 ;
        RECT 66.095 134.530 66.425 134.840 ;
        RECT 66.095 134.250 68.010 134.530 ;
        RECT 66.095 133.940 66.425 134.250 ;
        RECT 67.680 133.360 68.010 134.250 ;
        RECT 72.135 132.975 72.465 137.255 ;
        RECT 75.035 135.255 75.405 135.455 ;
        RECT 73.560 134.975 75.405 135.255 ;
        RECT 76.300 135.135 76.800 135.415 ;
        RECT 81.990 135.135 82.490 135.415 ;
        RECT 83.385 135.255 83.755 135.455 ;
        RECT 75.035 134.775 75.405 134.975 ;
        RECT 83.385 134.975 85.230 135.255 ;
        RECT 83.385 134.775 83.755 134.975 ;
        RECT 86.325 132.975 86.655 137.255 ;
        RECT 97.050 136.975 99.535 137.255 ;
        RECT 100.640 136.975 101.640 137.255 ;
        RECT 88.630 136.285 89.630 136.565 ;
        RECT 92.885 136.285 93.385 136.565 ;
        RECT 88.630 135.005 89.630 135.285 ;
        RECT 92.885 135.005 93.385 135.285 ;
        RECT 92.365 134.530 92.695 134.840 ;
        RECT 90.780 134.250 92.695 134.530 ;
        RECT 90.780 133.360 91.110 134.250 ;
        RECT 92.365 133.940 92.695 134.250 ;
        RECT 93.575 134.695 98.050 134.975 ;
        RECT 93.575 134.075 93.905 134.695 ;
        RECT 69.160 132.695 74.060 132.975 ;
        RECT 84.730 132.695 89.630 132.975 ;
        RECT 99.205 132.695 99.535 136.975 ;
        RECT 123.680 136.945 124.010 141.225 ;
        RECT 124.180 138.945 124.880 139.225 ;
        RECT 109.605 136.665 110.305 136.945 ;
        RECT 110.975 136.665 111.675 136.945 ;
        RECT 112.345 136.665 113.045 136.945 ;
        RECT 122.810 136.665 124.880 136.945 ;
        RECT 100.640 134.695 101.640 134.975 ;
        RECT 109.605 134.385 114.615 134.665 ;
        RECT 122.810 134.385 123.510 134.665 ;
        RECT 57.150 132.415 58.150 132.695 ;
        RECT 59.255 132.415 61.740 132.695 ;
        RECT 97.050 132.415 99.535 132.695 ;
        RECT 100.640 132.415 101.640 132.695 ;
        RECT 57.150 130.135 58.150 130.415 ;
        RECT 56.100 128.160 56.430 129.000 ;
        RECT 56.630 128.160 56.960 128.445 ;
        RECT 56.100 127.830 56.960 128.160 ;
        RECT 59.255 128.135 59.585 132.415 ;
        RECT 67.000 131.480 67.330 132.370 ;
        RECT 68.640 131.480 68.970 131.790 ;
        RECT 67.000 131.200 68.970 131.480 ;
        RECT 68.640 130.890 68.970 131.200 ;
        RECT 89.820 131.480 90.150 131.790 ;
        RECT 91.460 131.480 91.790 132.370 ;
        RECT 89.820 131.200 91.790 131.480 ;
        RECT 65.405 130.445 65.905 130.725 ;
        RECT 69.160 130.445 70.160 130.725 ;
        RECT 75.035 130.695 75.405 130.895 ;
        RECT 73.560 130.415 75.405 130.695 ;
        RECT 60.740 130.135 63.435 130.415 ;
        RECT 75.035 130.215 75.405 130.415 ;
        RECT 83.385 130.695 83.755 130.895 ;
        RECT 89.820 130.890 90.150 131.200 ;
        RECT 83.385 130.415 85.230 130.695 ;
        RECT 88.630 130.445 89.630 130.725 ;
        RECT 92.885 130.445 93.385 130.725 ;
        RECT 83.385 130.215 83.755 130.415 ;
        RECT 95.355 130.135 98.050 130.415 ;
        RECT 65.405 129.165 65.905 129.445 ;
        RECT 69.160 129.165 70.160 129.445 ;
        RECT 73.560 129.135 74.060 129.415 ;
        RECT 84.730 129.135 85.230 129.415 ;
        RECT 88.630 129.165 89.630 129.445 ;
        RECT 92.885 129.165 93.385 129.445 ;
        RECT 57.150 127.855 61.740 128.135 ;
        RECT 65.405 127.885 65.905 128.165 ;
        RECT 69.160 127.885 70.160 128.165 ;
        RECT 75.055 128.135 75.385 128.580 ;
        RECT 83.405 128.135 83.735 128.580 ;
        RECT 73.560 127.855 74.060 128.135 ;
        RECT 75.055 127.855 76.800 128.135 ;
        RECT 81.990 127.855 83.735 128.135 ;
        RECT 84.730 127.855 85.230 128.135 ;
        RECT 88.630 127.885 89.630 128.165 ;
        RECT 92.885 127.885 93.385 128.165 ;
        RECT 99.205 128.135 99.535 132.415 ;
        RECT 109.605 132.105 110.305 132.385 ;
        RECT 110.975 132.105 111.675 132.385 ;
        RECT 112.345 132.105 113.045 132.385 ;
        RECT 100.640 130.135 101.640 130.415 ;
        RECT 114.285 130.105 114.615 134.385 ;
        RECT 123.680 132.385 124.010 136.665 ;
        RECT 124.180 134.385 124.880 134.665 ;
        RECT 122.810 132.105 124.880 132.385 ;
        RECT 109.605 129.825 114.615 130.105 ;
        RECT 122.810 129.825 123.510 130.105 ;
        RECT 101.830 128.160 102.160 128.445 ;
        RECT 102.360 128.160 102.690 129.000 ;
        RECT 97.050 127.855 101.640 128.135 ;
        RECT 56.630 127.545 56.960 127.830 ;
        RECT 57.150 125.575 58.150 125.855 ;
        RECT 59.255 123.575 59.585 127.855 ;
        RECT 75.055 127.410 75.385 127.855 ;
        RECT 83.405 127.410 83.735 127.855 ;
        RECT 76.990 126.935 77.320 127.045 ;
        RECT 81.470 126.935 81.800 127.045 ;
        RECT 65.405 126.605 65.905 126.885 ;
        RECT 69.160 126.605 70.160 126.885 ;
        RECT 73.560 126.575 74.060 126.855 ;
        RECT 76.990 125.935 77.830 126.935 ;
        RECT 80.960 125.935 81.800 126.935 ;
        RECT 84.730 126.575 85.230 126.855 ;
        RECT 88.630 126.605 89.630 126.885 ;
        RECT 92.885 126.605 93.385 126.885 ;
        RECT 60.740 125.575 63.435 125.855 ;
        RECT 76.990 125.825 77.320 125.935 ;
        RECT 81.470 125.825 81.800 125.935 ;
        RECT 65.405 125.325 65.905 125.605 ;
        RECT 69.160 125.325 70.160 125.605 ;
        RECT 75.035 125.575 75.405 125.775 ;
        RECT 73.560 125.295 75.405 125.575 ;
        RECT 75.035 125.095 75.405 125.295 ;
        RECT 83.385 125.575 83.755 125.775 ;
        RECT 83.385 125.295 85.230 125.575 ;
        RECT 88.630 125.325 89.630 125.605 ;
        RECT 92.885 125.325 93.385 125.605 ;
        RECT 95.355 125.575 98.050 125.855 ;
        RECT 83.385 125.095 83.755 125.295 ;
        RECT 57.150 123.295 58.150 123.575 ;
        RECT 59.255 123.295 61.740 123.575 ;
        RECT 63.085 123.325 63.415 123.770 ;
        RECT 63.765 123.325 64.095 124.215 ;
        RECT 64.880 123.325 65.210 123.635 ;
        RECT 93.580 123.325 93.910 123.635 ;
        RECT 94.695 123.325 95.025 124.215 ;
        RECT 95.375 123.325 95.705 123.770 ;
        RECT 99.205 123.575 99.535 127.855 ;
        RECT 101.830 127.830 102.690 128.160 ;
        RECT 101.830 127.545 102.160 127.830 ;
        RECT 109.605 127.545 110.305 127.825 ;
        RECT 110.975 127.545 111.675 127.825 ;
        RECT 112.345 127.545 113.045 127.825 ;
        RECT 100.640 125.575 101.640 125.855 ;
        RECT 114.285 125.545 114.615 129.825 ;
        RECT 123.680 127.825 124.010 132.105 ;
        RECT 124.180 129.825 124.880 130.105 ;
        RECT 122.810 127.545 124.880 127.825 ;
        RECT 109.605 125.265 114.615 125.545 ;
        RECT 122.810 125.265 123.510 125.545 ;
        RECT 124.180 125.265 124.880 125.545 ;
        RECT 57.150 121.015 58.150 121.295 ;
        RECT 59.255 119.015 59.585 123.295 ;
        RECT 63.085 123.045 65.905 123.325 ;
        RECT 63.085 122.600 63.415 123.045 ;
        RECT 64.880 122.735 65.210 123.045 ;
        RECT 69.160 123.015 74.060 123.295 ;
        RECT 84.730 123.015 89.630 123.295 ;
        RECT 92.885 123.045 95.705 123.325 ;
        RECT 97.050 123.295 99.535 123.575 ;
        RECT 100.640 123.295 101.640 123.575 ;
        RECT 60.740 121.015 63.435 121.295 ;
        RECT 65.405 120.765 65.905 121.045 ;
        RECT 69.160 120.765 70.160 121.045 ;
        RECT 65.405 119.485 65.905 119.765 ;
        RECT 69.160 119.485 70.160 119.765 ;
        RECT 57.150 118.735 58.150 119.015 ;
        RECT 59.255 118.735 61.740 119.015 ;
        RECT 71.310 118.735 71.640 123.015 ;
        RECT 75.035 121.015 75.405 121.215 ;
        RECT 73.560 120.735 75.405 121.015 ;
        RECT 83.385 121.015 83.755 121.215 ;
        RECT 75.035 120.535 75.405 120.735 ;
        RECT 76.300 120.575 76.800 120.855 ;
        RECT 81.990 120.575 82.490 120.855 ;
        RECT 83.385 120.735 85.230 121.015 ;
        RECT 83.385 120.535 83.755 120.735 ;
        RECT 87.150 118.735 87.480 123.015 ;
        RECT 93.580 122.735 93.910 123.045 ;
        RECT 95.375 122.600 95.705 123.045 ;
        RECT 88.630 120.765 89.630 121.045 ;
        RECT 92.885 120.765 93.385 121.045 ;
        RECT 95.355 121.015 98.050 121.295 ;
        RECT 88.630 119.485 89.630 119.765 ;
        RECT 92.885 119.485 93.385 119.765 ;
        RECT 99.205 119.015 99.535 123.295 ;
        RECT 109.605 122.985 110.305 123.265 ;
        RECT 110.975 122.985 111.675 123.265 ;
        RECT 112.345 122.985 113.045 123.265 ;
        RECT 100.640 121.015 101.640 121.295 ;
        RECT 114.285 120.985 114.615 125.265 ;
        RECT 109.605 120.705 114.615 120.985 ;
        RECT 97.050 118.735 99.535 119.015 ;
        RECT 100.640 118.735 101.640 119.015 ;
        RECT 57.150 116.455 58.150 116.735 ;
        RECT 59.255 114.455 59.585 118.735 ;
        RECT 65.405 118.205 65.905 118.485 ;
        RECT 69.160 118.205 70.160 118.485 ;
        RECT 71.310 118.455 74.060 118.735 ;
        RECT 84.730 118.455 87.480 118.735 ;
        RECT 88.630 118.205 89.630 118.485 ;
        RECT 92.885 118.205 93.385 118.485 ;
        RECT 65.405 117.530 65.905 117.820 ;
        RECT 69.160 117.530 70.160 117.820 ;
        RECT 76.300 117.295 76.800 117.575 ;
        RECT 81.990 117.295 82.490 117.575 ;
        RECT 88.630 117.530 89.630 117.820 ;
        RECT 92.885 117.530 93.385 117.820 ;
        RECT 60.740 116.455 63.435 116.735 ;
        RECT 75.035 116.455 75.405 116.655 ;
        RECT 73.560 116.175 75.405 116.455 ;
        RECT 75.035 115.975 75.405 116.175 ;
        RECT 83.385 116.455 83.755 116.655 ;
        RECT 95.355 116.455 98.050 116.735 ;
        RECT 83.385 116.175 85.230 116.455 ;
        RECT 83.385 115.975 83.755 116.175 ;
        RECT 61.930 114.950 62.260 115.520 ;
        RECT 73.040 114.950 73.370 115.200 ;
        RECT 85.420 114.950 85.750 115.200 ;
        RECT 96.530 114.950 96.860 115.520 ;
        RECT 61.930 114.620 96.860 114.950 ;
        RECT 99.205 114.455 99.535 118.735 ;
        RECT 109.605 118.425 110.305 118.705 ;
        RECT 110.975 118.425 111.675 118.705 ;
        RECT 112.345 118.425 113.045 118.705 ;
        RECT 100.640 116.455 101.640 116.735 ;
        RECT 114.285 116.460 114.615 120.705 ;
        RECT 121.785 122.985 124.880 123.265 ;
        RECT 121.785 118.705 122.065 122.985 ;
        RECT 122.810 120.705 123.510 120.985 ;
        RECT 124.180 120.705 124.880 120.985 ;
        RECT 121.785 118.425 124.880 118.705 ;
        RECT 115.375 116.660 115.705 117.430 ;
        RECT 115.895 116.610 118.045 116.890 ;
        RECT 114.285 116.425 116.595 116.460 ;
        RECT 109.605 116.180 116.595 116.425 ;
        RECT 109.605 116.145 114.615 116.180 ;
        RECT 57.150 114.175 58.150 114.455 ;
        RECT 59.255 114.175 61.740 114.455 ;
        RECT 76.300 114.015 76.800 114.295 ;
        RECT 81.990 114.015 82.490 114.295 ;
        RECT 97.050 114.175 99.535 114.455 ;
        RECT 100.640 114.175 101.640 114.455 ;
        RECT 60.740 113.395 61.740 113.675 ;
        RECT 73.560 113.615 74.060 113.895 ;
        RECT 84.730 113.615 85.230 113.895 ;
        RECT 109.605 113.865 110.305 114.145 ;
        RECT 110.975 113.865 111.675 114.145 ;
        RECT 112.345 113.865 113.045 114.145 ;
        RECT 64.315 113.280 65.315 113.570 ;
        RECT 69.115 113.280 69.615 113.570 ;
        RECT 89.175 113.280 89.675 113.570 ;
        RECT 93.475 113.280 94.475 113.570 ;
        RECT 97.050 113.395 98.050 113.675 ;
        RECT 73.560 112.980 74.060 113.270 ;
        RECT 76.300 112.980 76.800 113.270 ;
        RECT 81.990 112.980 82.490 113.270 ;
        RECT 84.730 112.980 85.230 113.270 ;
        RECT 60.740 112.615 61.740 112.895 ;
        RECT 64.315 112.615 65.315 112.895 ;
        RECT 69.115 112.615 69.615 112.895 ;
        RECT 89.175 112.615 89.675 112.895 ;
        RECT 93.475 112.615 94.475 112.895 ;
        RECT 97.050 112.615 98.050 112.895 ;
        RECT 57.150 111.940 58.150 112.230 ;
        RECT 60.740 111.940 61.740 112.230 ;
        RECT 97.050 111.940 98.050 112.230 ;
        RECT 100.640 111.940 101.640 112.230 ;
        RECT 114.285 111.865 114.615 116.145 ;
        RECT 117.715 116.030 118.045 116.610 ;
        RECT 115.895 115.750 118.045 116.030 ;
        RECT 117.715 114.505 118.045 115.750 ;
        RECT 117.715 114.225 120.165 114.505 ;
        RECT 117.715 113.645 118.045 114.225 ;
        RECT 117.715 113.365 120.165 113.645 ;
        RECT 117.715 112.220 118.045 113.365 ;
        RECT 120.355 113.355 120.685 114.525 ;
        RECT 121.785 114.145 122.065 118.425 ;
        RECT 122.810 116.145 123.510 116.425 ;
        RECT 124.180 116.145 124.880 116.425 ;
        RECT 121.785 113.865 124.880 114.145 ;
        RECT 115.895 111.940 118.045 112.220 ;
        RECT 109.605 111.790 114.615 111.865 ;
        RECT 109.605 111.585 116.595 111.790 ;
        RECT 114.285 111.510 116.595 111.585 ;
        RECT 64.315 110.335 65.315 110.615 ;
        RECT 69.115 110.335 69.615 110.615 ;
        RECT 89.175 110.335 89.675 110.615 ;
        RECT 93.475 110.335 94.475 110.615 ;
        RECT 109.605 109.305 110.305 109.585 ;
        RECT 110.975 109.305 111.675 109.585 ;
        RECT 112.345 109.305 113.045 109.585 ;
        RECT 64.315 108.055 65.315 108.335 ;
        RECT 69.115 108.055 69.615 108.335 ;
        RECT 89.175 108.055 89.675 108.335 ;
        RECT 93.475 108.055 94.475 108.335 ;
        RECT 65.505 107.580 65.835 107.890 ;
        RECT 67.000 107.580 67.330 108.025 ;
        RECT 65.505 107.300 67.330 107.580 ;
        RECT 65.505 106.990 65.835 107.300 ;
        RECT 67.000 106.855 67.330 107.300 ;
        RECT 67.680 107.580 68.010 108.025 ;
        RECT 68.595 107.580 68.925 107.890 ;
        RECT 67.680 107.300 68.925 107.580 ;
        RECT 67.680 106.855 68.010 107.300 ;
        RECT 68.595 106.990 68.925 107.300 ;
        RECT 89.865 107.580 90.195 107.890 ;
        RECT 90.780 107.580 91.110 108.025 ;
        RECT 89.865 107.300 91.110 107.580 ;
        RECT 89.865 106.990 90.195 107.300 ;
        RECT 90.780 106.855 91.110 107.300 ;
        RECT 91.460 107.580 91.790 108.025 ;
        RECT 92.955 107.580 93.285 107.890 ;
        RECT 91.460 107.300 93.285 107.580 ;
        RECT 114.285 107.305 114.615 111.510 ;
        RECT 117.715 111.360 118.045 111.940 ;
        RECT 115.895 111.080 118.045 111.360 ;
        RECT 116.785 110.110 117.115 110.880 ;
        RECT 91.460 106.855 91.790 107.300 ;
        RECT 92.955 106.990 93.285 107.300 ;
        RECT 109.605 107.025 114.615 107.305 ;
        RECT 64.315 105.775 69.615 106.055 ;
        RECT 89.175 105.775 94.475 106.055 ;
        RECT 109.605 104.745 110.305 105.025 ;
        RECT 110.975 104.745 111.675 105.025 ;
        RECT 112.345 104.745 113.045 105.025 ;
        RECT 64.315 103.495 65.315 103.775 ;
        RECT 69.115 103.495 69.615 103.775 ;
        RECT 89.175 103.495 89.675 103.775 ;
        RECT 93.475 103.495 94.475 103.775 ;
        RECT 114.285 102.745 114.615 107.025 ;
        RECT 109.605 102.465 114.615 102.745 ;
        RECT 64.315 101.215 69.615 101.495 ;
        RECT 89.175 101.215 94.475 101.495 ;
        RECT 109.605 100.185 110.305 100.465 ;
        RECT 110.975 100.185 111.675 100.465 ;
        RECT 112.345 100.185 113.045 100.465 ;
        RECT 114.285 100.090 114.615 102.465 ;
        RECT 121.785 109.585 122.065 113.865 ;
        RECT 122.810 111.585 123.510 111.865 ;
        RECT 124.180 111.585 124.880 111.865 ;
        RECT 121.785 109.305 124.880 109.585 ;
        RECT 121.785 105.025 122.065 109.305 ;
        RECT 122.810 107.025 123.510 107.305 ;
        RECT 124.180 107.025 124.880 107.305 ;
        RECT 121.785 104.745 124.880 105.025 ;
        RECT 121.785 100.465 122.065 104.745 ;
        RECT 122.810 102.465 123.510 102.745 ;
        RECT 124.180 102.465 124.880 102.745 ;
        RECT 121.785 100.185 124.880 100.465 ;
        RECT 111.845 99.395 112.175 99.755 ;
        RECT 121.785 99.395 122.065 100.185 ;
        RECT 64.315 98.935 65.315 99.215 ;
        RECT 69.115 98.935 69.615 99.215 ;
        RECT 89.175 98.935 89.675 99.215 ;
        RECT 93.475 98.935 94.475 99.215 ;
        RECT 111.845 98.895 122.065 99.395 ;
        RECT 111.845 98.535 112.175 98.895 ;
        RECT 109.605 97.905 114.615 98.185 ;
        RECT 64.315 96.655 69.615 96.935 ;
        RECT 89.175 96.655 94.475 96.935 ;
        RECT 109.605 95.625 110.305 95.905 ;
        RECT 110.975 95.625 111.675 95.905 ;
        RECT 112.345 95.625 113.045 95.905 ;
        RECT 64.315 94.375 65.315 94.655 ;
        RECT 69.115 94.375 69.615 94.655 ;
        RECT 89.175 94.375 89.675 94.655 ;
        RECT 93.475 94.375 94.475 94.655 ;
        RECT 114.285 93.625 114.615 97.905 ;
        RECT 109.605 93.345 114.615 93.625 ;
        RECT 121.785 95.905 122.065 98.895 ;
        RECT 122.810 97.905 123.510 98.185 ;
        RECT 124.180 97.905 124.880 98.185 ;
        RECT 121.785 95.625 124.880 95.905 ;
        RECT 64.315 92.095 65.315 92.375 ;
        RECT 69.115 92.095 69.615 92.375 ;
        RECT 89.175 92.095 89.675 92.375 ;
        RECT 93.475 92.095 94.475 92.375 ;
        RECT 121.785 91.345 122.065 95.625 ;
        RECT 122.810 93.345 123.510 93.625 ;
        RECT 124.180 93.345 124.880 93.625 ;
        RECT 109.605 91.065 110.305 91.345 ;
        RECT 110.975 91.065 111.675 91.345 ;
        RECT 112.345 91.065 113.045 91.345 ;
        RECT 121.785 91.065 124.880 91.345 ;
        RECT 64.315 89.815 65.315 90.095 ;
        RECT 69.115 89.815 69.615 90.095 ;
        RECT 89.175 89.815 89.675 90.095 ;
        RECT 93.475 89.815 94.475 90.095 ;
        RECT 64.315 89.140 65.315 89.430 ;
        RECT 69.115 89.140 69.615 89.430 ;
        RECT 89.175 89.140 89.675 89.430 ;
        RECT 93.475 89.140 94.475 89.430 ;
        RECT 109.605 88.785 114.615 89.065 ;
        RECT 122.810 88.785 123.510 89.065 ;
        RECT 124.180 88.785 124.880 89.065 ;
        RECT 79.165 86.490 104.670 87.090 ;
        RECT 109.605 86.505 110.305 86.785 ;
        RECT 110.975 86.505 111.675 86.785 ;
        RECT 112.345 86.505 113.045 86.785 ;
        RECT 104.070 86.010 104.670 86.490 ;
        RECT 83.780 84.955 88.005 85.285 ;
        RECT 74.410 83.825 87.435 84.155 ;
        RECT 71.925 83.245 78.995 83.525 ;
        RECT 79.565 83.245 86.635 83.525 ;
        RECT 71.925 82.355 72.255 83.245 ;
        RECT 72.595 82.610 73.445 82.900 ;
        RECT 75.820 82.610 76.670 82.900 ;
        RECT 77.395 82.610 78.245 82.900 ;
        RECT 78.585 82.355 78.915 83.245 ;
        RECT 79.645 82.355 79.975 83.245 ;
        RECT 80.315 82.610 81.165 82.900 ;
        RECT 81.890 82.610 82.740 82.900 ;
        RECT 85.115 82.610 85.965 82.900 ;
        RECT 86.305 82.355 86.635 83.245 ;
        RECT 72.595 81.945 73.445 82.225 ;
        RECT 72.595 81.515 73.445 81.795 ;
        RECT 71.905 80.455 72.275 81.135 ;
        RECT 72.595 81.085 73.445 81.365 ;
        RECT 74.430 81.285 74.760 82.145 ;
        RECT 75.820 81.945 76.670 82.225 ;
        RECT 77.395 81.945 78.245 82.225 ;
        RECT 80.315 81.945 81.165 82.225 ;
        RECT 81.890 81.945 82.740 82.225 ;
        RECT 75.820 81.515 76.670 81.795 ;
        RECT 77.395 81.515 78.245 81.795 ;
        RECT 80.315 81.515 81.165 81.795 ;
        RECT 81.890 81.515 82.740 81.795 ;
        RECT 75.745 81.085 77.215 81.365 ;
        RECT 77.395 81.085 78.245 81.365 ;
        RECT 76.925 80.935 77.215 81.085 ;
        RECT 72.445 80.655 76.745 80.935 ;
        RECT 76.925 80.655 78.395 80.935 ;
        RECT 72.595 80.225 73.445 80.505 ;
        RECT 74.430 80.075 74.760 80.655 ;
        RECT 76.925 80.505 77.215 80.655 ;
        RECT 75.745 80.225 77.215 80.505 ;
        RECT 77.395 80.225 78.245 80.505 ;
        RECT 76.925 80.075 77.215 80.225 ;
        RECT 72.445 79.795 76.745 80.075 ;
        RECT 76.925 79.795 78.395 80.075 ;
        RECT 72.595 79.365 73.445 79.645 ;
        RECT 72.595 78.935 73.445 79.215 ;
        RECT 72.595 78.505 73.445 78.785 ;
        RECT 72.595 77.830 73.445 78.135 ;
        RECT 74.430 77.685 74.760 79.795 ;
        RECT 76.925 79.645 77.215 79.795 ;
        RECT 75.745 79.365 77.215 79.645 ;
        RECT 77.395 79.365 78.245 79.645 ;
        RECT 78.585 79.640 78.915 81.090 ;
        RECT 79.645 79.640 79.975 81.090 ;
        RECT 80.315 81.085 81.165 81.365 ;
        RECT 81.345 81.085 82.815 81.365 ;
        RECT 83.800 81.285 84.130 82.145 ;
        RECT 85.115 81.945 85.965 82.225 ;
        RECT 85.115 81.515 85.965 81.795 ;
        RECT 85.115 81.085 85.965 81.365 ;
        RECT 81.345 80.935 81.635 81.085 ;
        RECT 80.165 80.655 81.635 80.935 ;
        RECT 81.815 80.655 86.115 80.935 ;
        RECT 81.345 80.505 81.635 80.655 ;
        RECT 80.315 80.225 81.165 80.505 ;
        RECT 81.345 80.225 82.815 80.505 ;
        RECT 81.345 80.075 81.635 80.225 ;
        RECT 83.800 80.075 84.130 80.655 ;
        RECT 85.115 80.225 85.965 80.505 ;
        RECT 86.285 80.455 86.655 81.135 ;
        RECT 80.165 79.795 81.635 80.075 ;
        RECT 81.815 79.795 86.115 80.075 ;
        RECT 81.345 79.645 81.635 79.795 ;
        RECT 80.315 79.365 81.165 79.645 ;
        RECT 81.345 79.365 82.815 79.645 ;
        RECT 75.820 78.935 76.670 79.215 ;
        RECT 77.395 78.935 78.245 79.215 ;
        RECT 80.315 78.935 81.165 79.215 ;
        RECT 81.890 78.935 82.740 79.215 ;
        RECT 75.820 78.505 76.670 78.785 ;
        RECT 77.395 78.505 78.245 78.785 ;
        RECT 80.315 78.505 81.165 78.785 ;
        RECT 81.890 78.505 82.740 78.785 ;
        RECT 75.820 77.830 76.670 78.135 ;
        RECT 77.395 77.830 78.245 78.135 ;
        RECT 80.315 77.830 81.165 78.135 ;
        RECT 81.890 77.830 82.740 78.135 ;
        RECT 83.800 77.685 84.130 79.795 ;
        RECT 85.115 79.365 85.965 79.645 ;
        RECT 85.115 78.935 85.965 79.215 ;
        RECT 85.115 78.505 85.965 78.785 ;
        RECT 85.115 77.830 85.965 78.135 ;
        RECT 87.085 77.685 87.415 78.525 ;
        RECT 74.430 77.355 79.995 77.685 ;
        RECT 83.800 77.355 87.415 77.685 ;
        RECT 76.360 75.680 76.690 77.355 ;
        RECT 87.675 77.240 88.005 84.955 ;
        RECT 114.285 84.505 114.615 88.785 ;
        RECT 122.810 86.505 123.510 86.785 ;
        RECT 124.180 86.505 124.880 86.785 ;
        RECT 109.605 84.225 114.615 84.505 ;
        RECT 122.810 84.225 123.510 84.505 ;
        RECT 124.180 84.225 124.880 84.505 ;
        RECT 89.110 82.960 90.110 83.250 ;
        RECT 92.960 82.960 93.960 83.250 ;
        RECT 89.110 82.295 90.110 82.575 ;
        RECT 89.110 81.865 90.110 82.145 ;
        RECT 91.120 81.795 91.450 82.565 ;
        RECT 92.960 82.295 93.960 82.575 ;
        RECT 114.285 82.260 114.615 84.225 ;
        RECT 122.330 83.360 122.620 83.700 ;
        RECT 123.680 83.360 124.010 83.670 ;
        RECT 115.375 82.460 115.705 83.230 ;
        RECT 122.330 83.080 124.010 83.360 ;
        RECT 122.330 82.740 122.620 83.080 ;
        RECT 123.680 82.770 124.010 83.080 ;
        RECT 115.895 82.410 118.045 82.690 ;
        RECT 92.960 81.865 93.960 82.145 ;
        RECT 109.605 81.945 110.305 82.225 ;
        RECT 110.975 81.945 111.675 82.225 ;
        RECT 112.345 81.945 113.045 82.225 ;
        RECT 114.285 81.980 116.595 82.260 ;
        RECT 89.110 81.435 90.110 81.715 ;
        RECT 92.960 81.435 93.960 81.715 ;
        RECT 89.110 81.005 94.460 81.285 ;
        RECT 89.110 80.575 90.110 80.855 ;
        RECT 91.120 80.425 91.450 81.005 ;
        RECT 92.960 80.575 93.960 80.855 ;
        RECT 89.110 80.145 94.460 80.425 ;
        RECT 89.110 79.715 90.110 79.995 ;
        RECT 89.110 79.285 90.110 79.565 ;
        RECT 89.110 78.855 90.110 79.135 ;
        RECT 89.110 78.180 90.110 78.470 ;
        RECT 91.120 77.240 91.450 80.145 ;
        RECT 92.960 79.715 93.960 79.995 ;
        RECT 114.285 79.945 114.615 81.980 ;
        RECT 117.715 81.830 118.045 82.410 ;
        RECT 115.895 81.550 118.045 81.830 ;
        RECT 109.605 79.665 114.615 79.945 ;
        RECT 92.960 79.285 93.960 79.565 ;
        RECT 92.960 78.855 93.960 79.135 ;
        RECT 92.960 78.180 93.960 78.470 ;
        RECT 109.605 77.385 110.305 77.665 ;
        RECT 110.975 77.385 111.675 77.665 ;
        RECT 112.345 77.385 113.045 77.665 ;
        RECT 114.285 77.590 114.615 79.665 ;
        RECT 117.715 80.305 118.045 81.550 ;
        RECT 121.155 81.945 123.510 82.225 ;
        RECT 124.180 81.945 124.880 82.225 ;
        RECT 121.155 81.055 121.485 81.945 ;
        RECT 117.715 80.025 120.165 80.305 ;
        RECT 117.715 79.445 118.045 80.025 ;
        RECT 117.715 79.165 120.165 79.445 ;
        RECT 117.715 78.020 118.045 79.165 ;
        RECT 120.355 79.155 120.685 80.325 ;
        RECT 122.810 79.665 123.510 79.945 ;
        RECT 124.180 79.665 124.880 79.945 ;
        RECT 115.895 77.740 118.045 78.020 ;
        RECT 87.675 76.910 91.450 77.240 ;
        RECT 114.285 77.310 116.595 77.590 ;
        RECT 91.120 75.095 95.795 75.425 ;
        RECT 114.285 75.385 114.615 77.310 ;
        RECT 117.715 77.160 118.045 77.740 ;
        RECT 122.810 77.385 123.510 77.665 ;
        RECT 124.180 77.385 124.880 77.665 ;
        RECT 115.895 76.880 118.045 77.160 ;
        RECT 122.810 76.750 123.510 77.040 ;
        RECT 124.180 76.750 124.880 77.040 ;
        RECT 116.785 75.910 117.115 76.680 ;
        RECT 109.605 75.105 114.615 75.385 ;
        RECT 115.745 75.345 116.445 75.635 ;
        RECT 91.120 74.255 91.450 75.095 ;
        RECT 109.605 72.825 110.305 73.105 ;
        RECT 110.975 72.825 111.675 73.105 ;
        RECT 112.345 72.825 113.045 73.105 ;
        RECT 65.330 72.300 66.330 72.590 ;
        RECT 69.180 72.300 70.180 72.590 ;
        RECT 74.350 72.300 75.350 72.590 ;
        RECT 78.200 72.300 79.200 72.590 ;
        RECT 81.290 72.300 82.290 72.590 ;
        RECT 85.140 72.300 86.140 72.590 ;
        RECT 89.110 72.300 90.110 72.590 ;
        RECT 92.960 72.300 93.960 72.590 ;
        RECT 65.330 71.635 66.330 71.915 ;
        RECT 65.330 71.205 66.330 71.485 ;
        RECT 67.340 71.135 67.670 71.905 ;
        RECT 69.180 71.635 70.180 71.915 ;
        RECT 74.350 71.635 75.350 71.915 ;
        RECT 69.180 71.205 70.180 71.485 ;
        RECT 74.350 71.205 75.350 71.485 ;
        RECT 76.360 71.135 76.690 71.905 ;
        RECT 78.200 71.635 79.200 71.915 ;
        RECT 81.290 71.635 82.290 71.915 ;
        RECT 78.200 71.205 79.200 71.485 ;
        RECT 81.290 71.205 82.290 71.485 ;
        RECT 83.800 71.135 84.130 71.905 ;
        RECT 85.140 71.635 86.140 71.915 ;
        RECT 89.110 71.635 90.110 71.915 ;
        RECT 85.140 71.205 86.140 71.485 ;
        RECT 89.110 71.205 90.110 71.485 ;
        RECT 91.120 71.135 91.450 71.905 ;
        RECT 92.960 71.635 93.960 71.915 ;
        RECT 92.960 71.205 93.960 71.485 ;
        RECT 65.330 70.775 66.330 71.055 ;
        RECT 69.180 70.775 70.180 71.055 ;
        RECT 74.350 70.775 75.350 71.055 ;
        RECT 78.200 70.775 79.200 71.055 ;
        RECT 81.290 70.775 82.290 71.055 ;
        RECT 85.140 70.775 86.140 71.055 ;
        RECT 89.110 70.775 90.110 71.055 ;
        RECT 92.960 70.775 93.960 71.055 ;
        RECT 114.285 70.825 114.615 75.105 ;
        RECT 120.330 71.200 124.290 71.530 ;
        RECT 65.330 70.345 70.680 70.625 ;
        RECT 74.350 70.345 79.700 70.625 ;
        RECT 80.790 70.345 86.140 70.625 ;
        RECT 89.110 70.345 94.460 70.625 ;
        RECT 109.605 70.545 114.615 70.825 ;
        RECT 115.745 70.570 116.445 70.860 ;
        RECT 65.330 69.915 66.330 70.195 ;
        RECT 67.340 69.765 67.670 70.345 ;
        RECT 69.180 69.915 70.180 70.195 ;
        RECT 74.350 69.915 75.350 70.195 ;
        RECT 76.360 69.765 76.690 70.345 ;
        RECT 78.200 69.915 79.200 70.195 ;
        RECT 81.290 69.915 82.290 70.195 ;
        RECT 83.800 69.765 84.130 70.345 ;
        RECT 85.140 69.915 86.140 70.195 ;
        RECT 89.110 69.915 90.110 70.195 ;
        RECT 91.120 69.765 91.450 70.345 ;
        RECT 119.440 70.290 120.140 70.580 ;
        RECT 92.960 69.915 93.960 70.195 ;
        RECT 65.330 69.485 70.680 69.765 ;
        RECT 74.350 69.485 79.700 69.765 ;
        RECT 80.790 69.485 86.140 69.765 ;
        RECT 89.110 69.485 94.460 69.765 ;
        RECT 111.845 69.690 112.175 70.000 ;
        RECT 115.745 69.905 116.445 70.185 ;
        RECT 111.845 69.410 115.555 69.690 ;
        RECT 119.440 69.625 120.140 69.905 ;
        RECT 65.330 69.055 66.330 69.335 ;
        RECT 69.180 69.055 70.180 69.335 ;
        RECT 74.350 69.055 75.350 69.335 ;
        RECT 78.200 69.055 79.200 69.335 ;
        RECT 81.290 69.055 82.290 69.335 ;
        RECT 85.140 69.055 86.140 69.335 ;
        RECT 89.110 69.055 90.110 69.335 ;
        RECT 92.960 69.055 93.960 69.335 ;
        RECT 111.845 69.100 112.175 69.410 ;
        RECT 65.330 68.625 70.680 68.905 ;
        RECT 74.350 68.625 79.700 68.905 ;
        RECT 80.790 68.625 86.140 68.905 ;
        RECT 89.110 68.625 94.460 68.905 ;
        RECT 115.225 68.790 115.555 69.410 ;
        RECT 119.440 69.195 120.140 69.475 ;
        RECT 120.330 69.400 120.660 71.200 ;
        RECT 123.960 70.360 124.290 71.200 ;
        RECT 125.425 70.250 126.125 70.540 ;
        RECT 117.715 68.765 120.140 69.045 ;
        RECT 121.155 68.765 122.855 69.045 ;
        RECT 123.045 69.020 123.375 70.055 ;
        RECT 125.425 69.625 126.125 69.905 ;
        RECT 125.425 69.195 126.125 69.475 ;
        RECT 125.425 68.765 126.125 69.045 ;
        RECT 65.330 68.195 66.330 68.475 ;
        RECT 67.340 68.045 67.670 68.625 ;
        RECT 69.180 68.195 70.180 68.475 ;
        RECT 74.350 68.195 75.350 68.475 ;
        RECT 76.360 68.045 76.690 68.625 ;
        RECT 78.200 68.195 79.200 68.475 ;
        RECT 81.290 68.195 82.290 68.475 ;
        RECT 83.800 68.045 84.130 68.625 ;
        RECT 85.140 68.195 86.140 68.475 ;
        RECT 89.110 68.195 90.110 68.475 ;
        RECT 91.120 68.045 91.450 68.625 ;
        RECT 92.960 68.195 93.960 68.475 ;
        RECT 109.605 68.265 110.305 68.545 ;
        RECT 110.975 68.265 111.675 68.545 ;
        RECT 112.345 68.265 113.045 68.545 ;
        RECT 117.715 68.185 118.045 68.765 ;
        RECT 119.440 68.615 120.140 68.620 ;
        RECT 119.440 68.335 124.290 68.615 ;
        RECT 125.425 68.335 126.125 68.615 ;
        RECT 65.330 67.765 70.680 68.045 ;
        RECT 74.350 67.765 79.700 68.045 ;
        RECT 80.790 67.765 86.140 68.045 ;
        RECT 89.110 67.765 94.460 68.045 ;
        RECT 117.715 67.905 120.140 68.185 ;
        RECT 121.155 67.905 122.855 68.185 ;
        RECT 65.330 67.335 66.330 67.615 ;
        RECT 67.340 67.185 67.670 67.765 ;
        RECT 69.180 67.335 70.180 67.615 ;
        RECT 74.350 67.335 75.350 67.615 ;
        RECT 76.360 67.185 76.690 67.765 ;
        RECT 78.200 67.335 79.200 67.615 ;
        RECT 81.290 67.335 82.290 67.615 ;
        RECT 83.800 67.185 84.130 67.765 ;
        RECT 85.140 67.335 86.140 67.615 ;
        RECT 89.110 67.335 90.110 67.615 ;
        RECT 91.120 67.185 91.450 67.765 ;
        RECT 115.745 67.625 116.445 67.905 ;
        RECT 92.960 67.335 93.960 67.615 ;
        RECT 117.715 67.325 118.045 67.905 ;
        RECT 119.440 67.755 120.140 67.760 ;
        RECT 123.960 67.755 124.290 68.335 ;
        RECT 125.425 67.905 126.125 68.185 ;
        RECT 119.440 67.475 124.290 67.755 ;
        RECT 125.425 67.475 126.125 67.755 ;
        RECT 65.330 66.905 70.680 67.185 ;
        RECT 74.350 66.905 79.700 67.185 ;
        RECT 80.790 66.905 86.140 67.185 ;
        RECT 89.110 66.905 94.460 67.185 ;
        RECT 117.715 67.045 120.140 67.325 ;
        RECT 121.155 67.045 122.855 67.325 ;
        RECT 65.330 66.475 66.330 66.755 ;
        RECT 67.340 66.325 67.670 66.905 ;
        RECT 69.180 66.475 70.180 66.755 ;
        RECT 74.350 66.475 75.350 66.755 ;
        RECT 76.360 66.325 76.690 66.905 ;
        RECT 78.200 66.475 79.200 66.755 ;
        RECT 81.290 66.475 82.290 66.755 ;
        RECT 83.800 66.325 84.130 66.905 ;
        RECT 85.140 66.475 86.140 66.755 ;
        RECT 89.110 66.475 90.110 66.755 ;
        RECT 91.120 66.325 91.450 66.905 ;
        RECT 92.960 66.475 93.960 66.755 ;
        RECT 65.330 66.045 70.680 66.325 ;
        RECT 74.350 66.045 79.700 66.325 ;
        RECT 80.790 66.045 86.140 66.325 ;
        RECT 89.110 66.045 94.460 66.325 ;
        RECT 65.330 65.615 66.330 65.895 ;
        RECT 67.340 65.465 67.670 66.045 ;
        RECT 69.180 65.615 70.180 65.895 ;
        RECT 74.350 65.615 75.350 65.895 ;
        RECT 76.360 65.465 76.690 66.045 ;
        RECT 78.200 65.615 79.200 65.895 ;
        RECT 81.290 65.615 82.290 65.895 ;
        RECT 83.800 65.465 84.130 66.045 ;
        RECT 85.140 65.615 86.140 65.895 ;
        RECT 89.110 65.615 90.110 65.895 ;
        RECT 91.120 65.465 91.450 66.045 ;
        RECT 109.605 65.985 110.305 66.265 ;
        RECT 110.975 65.985 111.675 66.265 ;
        RECT 112.345 65.985 113.045 66.265 ;
        RECT 92.960 65.615 93.960 65.895 ;
        RECT 117.715 65.625 118.045 67.045 ;
        RECT 119.440 66.615 120.140 66.895 ;
        RECT 119.440 66.185 120.140 66.465 ;
        RECT 65.330 65.185 70.680 65.465 ;
        RECT 74.350 65.185 79.700 65.465 ;
        RECT 80.790 65.185 86.140 65.465 ;
        RECT 89.110 65.185 94.460 65.465 ;
        RECT 115.745 65.345 118.045 65.625 ;
        RECT 65.330 64.755 66.330 65.035 ;
        RECT 65.330 64.325 66.330 64.605 ;
        RECT 65.330 63.895 66.330 64.175 ;
        RECT 67.340 63.950 67.670 65.185 ;
        RECT 69.180 64.755 70.180 65.035 ;
        RECT 74.350 64.755 75.350 65.035 ;
        RECT 69.180 64.325 70.180 64.605 ;
        RECT 74.350 64.325 75.350 64.605 ;
        RECT 69.180 63.895 70.180 64.175 ;
        RECT 74.350 63.895 75.350 64.175 ;
        RECT 76.360 63.950 76.690 65.185 ;
        RECT 78.200 64.755 79.200 65.035 ;
        RECT 81.290 64.755 82.290 65.035 ;
        RECT 78.200 64.325 79.200 64.605 ;
        RECT 81.290 64.325 82.290 64.605 ;
        RECT 78.200 63.895 79.200 64.175 ;
        RECT 81.290 63.895 82.290 64.175 ;
        RECT 83.800 63.950 84.130 65.185 ;
        RECT 85.140 64.755 86.140 65.035 ;
        RECT 89.110 64.755 90.110 65.035 ;
        RECT 85.140 64.325 86.140 64.605 ;
        RECT 89.110 64.325 90.110 64.605 ;
        RECT 85.140 63.895 86.140 64.175 ;
        RECT 89.110 63.895 90.110 64.175 ;
        RECT 91.120 63.950 91.450 65.185 ;
        RECT 92.960 64.755 93.960 65.035 ;
        RECT 92.960 64.325 93.960 64.605 ;
        RECT 92.960 63.895 93.960 64.175 ;
        RECT 109.605 63.705 110.305 63.985 ;
        RECT 110.975 63.705 111.675 63.985 ;
        RECT 112.345 63.705 113.045 63.985 ;
        RECT 117.715 63.795 118.045 65.345 ;
        RECT 123.960 66.035 124.290 67.475 ;
        RECT 125.425 67.045 126.125 67.325 ;
        RECT 125.425 66.615 126.125 66.895 ;
        RECT 125.425 66.185 126.125 66.465 ;
        RECT 123.960 65.755 126.125 66.035 ;
        RECT 123.960 65.175 124.290 65.755 ;
        RECT 124.640 65.175 125.240 65.755 ;
        RECT 126.305 65.615 126.625 65.900 ;
        RECT 127.395 65.615 127.725 66.035 ;
        RECT 125.425 65.325 126.125 65.605 ;
        RECT 126.305 65.285 127.725 65.615 ;
        RECT 123.960 64.895 126.125 65.175 ;
        RECT 126.305 65.000 126.625 65.285 ;
        RECT 119.440 64.375 120.140 64.655 ;
        RECT 119.440 63.945 120.140 64.225 ;
        RECT 117.715 63.515 120.140 63.795 ;
        RECT 120.440 63.625 120.770 64.715 ;
        RECT 121.155 63.515 122.855 63.795 ;
        RECT 65.330 63.220 66.330 63.510 ;
        RECT 69.180 63.220 70.180 63.510 ;
        RECT 74.350 63.220 75.350 63.510 ;
        RECT 78.200 63.220 79.200 63.510 ;
        RECT 81.290 63.220 82.290 63.510 ;
        RECT 85.140 63.220 86.140 63.510 ;
        RECT 89.110 63.220 90.110 63.510 ;
        RECT 92.960 63.220 93.960 63.510 ;
        RECT 109.605 63.030 110.305 63.320 ;
        RECT 110.975 63.030 111.675 63.320 ;
        RECT 112.345 63.030 113.045 63.320 ;
        RECT 115.745 63.065 116.445 63.345 ;
        RECT 117.715 62.935 118.045 63.515 ;
        RECT 119.440 63.365 120.140 63.370 ;
        RECT 123.960 63.365 124.290 64.895 ;
        RECT 119.440 63.085 124.290 63.365 ;
        RECT 117.715 62.655 120.140 62.935 ;
        RECT 121.155 62.655 122.855 62.935 ;
        RECT 117.715 62.075 118.045 62.655 ;
        RECT 119.440 62.505 120.140 62.510 ;
        RECT 123.960 62.505 124.290 63.085 ;
        RECT 119.440 62.225 124.290 62.505 ;
        RECT 117.715 61.795 120.140 62.075 ;
        RECT 121.135 61.795 122.855 62.075 ;
        RECT 119.440 61.365 120.140 61.645 ;
        RECT 123.045 61.555 123.375 61.680 ;
        RECT 123.940 61.555 124.310 61.730 ;
        RECT 123.045 61.225 124.310 61.555 ;
        RECT 115.745 60.785 116.445 61.065 ;
        RECT 119.440 60.935 120.140 61.215 ;
        RECT 123.045 61.100 123.375 61.225 ;
        RECT 123.940 61.050 124.310 61.225 ;
        RECT 115.745 60.110 116.445 60.400 ;
        RECT 119.440 60.300 120.140 60.590 ;
        RECT 120.420 59.400 123.395 59.730 ;
        RECT 124.640 55.515 125.240 64.895 ;
        RECT 127.395 64.865 127.725 65.285 ;
        RECT 125.425 64.465 126.125 64.745 ;
        RECT 125.425 64.035 126.125 64.315 ;
        RECT 125.425 63.605 126.125 63.885 ;
        RECT 125.425 63.175 126.125 63.455 ;
        RECT 125.425 62.745 126.125 63.025 ;
        RECT 125.425 62.315 126.125 62.595 ;
        RECT 125.425 61.885 126.125 62.165 ;
        RECT 125.425 61.455 126.125 61.735 ;
        RECT 125.425 61.025 126.125 61.305 ;
        RECT 125.425 60.390 126.125 60.680 ;
        RECT 124.640 38.705 142.530 39.305 ;
        RECT 104.070 21.455 104.670 21.960 ;
        RECT 124.640 21.455 125.240 21.695 ;
        RECT 72.280 20.305 72.610 21.145 ;
        RECT 104.070 20.855 125.240 21.455 ;
        RECT 124.640 20.615 125.240 20.855 ;
        RECT 72.280 19.975 124.290 20.305 ;
        RECT 87.515 19.145 123.375 19.475 ;
        RECT 123.960 19.135 124.290 19.975 ;
        RECT 105.170 18.045 118.045 18.645 ;
        RECT 90.985 16.475 91.585 16.955 ;
        RECT 47.095 15.875 91.585 16.475 ;
        RECT 45.995 14.775 84.265 15.375 ;
        RECT 117.715 13.545 142.530 14.145 ;
        RECT 76.225 7.495 113.000 8.095 ;
        RECT 67.205 6.395 90.920 6.995 ;
        RECT 157.665 4.675 158.265 5.555 ;
        RECT 134.480 4.075 158.265 4.675 ;
      LAYER via2 ;
        RECT 127.420 211.825 127.700 212.105 ;
        RECT 127.820 211.825 128.100 212.105 ;
        RECT 128.220 211.825 128.500 212.105 ;
        RECT 143.030 211.825 143.310 212.105 ;
        RECT 143.430 211.825 143.710 212.105 ;
        RECT 143.830 211.825 144.110 212.105 ;
        RECT 115.400 210.995 115.680 211.275 ;
        RECT 115.800 210.995 116.080 211.275 ;
        RECT 116.200 210.995 116.480 211.275 ;
        RECT 157.825 211.020 158.105 211.300 ;
        RECT 157.825 210.620 158.105 210.900 ;
        RECT 120.380 210.165 120.660 210.445 ;
        RECT 120.780 210.165 121.060 210.445 ;
        RECT 121.180 210.165 121.460 210.445 ;
        RECT 146.705 210.165 146.985 210.445 ;
        RECT 147.105 210.165 147.385 210.445 ;
        RECT 147.505 210.165 147.785 210.445 ;
        RECT 157.825 210.220 158.105 210.500 ;
        RECT 123.705 209.200 123.985 209.480 ;
        RECT 124.105 209.200 124.385 209.480 ;
        RECT 156.725 209.360 157.005 209.640 ;
        RECT 156.725 208.960 157.005 209.240 ;
        RECT 117.740 208.100 118.020 208.380 ;
        RECT 118.140 208.100 118.420 208.380 ;
        RECT 118.540 208.100 118.820 208.380 ;
        RECT 140.825 208.100 141.105 208.380 ;
        RECT 141.225 208.100 141.505 208.380 ;
        RECT 141.625 208.100 141.905 208.380 ;
        RECT 142.025 208.100 142.305 208.380 ;
        RECT 106.125 206.605 106.405 206.885 ;
        RECT 106.525 206.605 106.805 206.885 ;
        RECT 106.925 206.605 107.205 206.885 ;
        RECT 117.740 206.765 118.020 207.045 ;
        RECT 117.740 206.365 118.020 206.645 ;
        RECT 117.740 205.965 118.020 206.245 ;
        RECT 84.960 174.565 85.240 174.845 ;
        RECT 84.960 174.165 85.240 174.445 ;
        RECT 84.960 173.765 85.240 174.045 ;
        RECT 108.355 173.845 108.635 174.125 ;
        RECT 108.755 173.845 109.035 174.125 ;
        RECT 112.205 173.845 112.485 174.125 ;
        RECT 112.605 173.845 112.885 174.125 ;
        RECT 88.640 173.465 88.920 173.745 ;
        RECT 88.640 173.065 88.920 173.345 ;
        RECT 108.355 173.175 108.635 173.455 ;
        RECT 108.755 173.175 109.035 173.455 ;
        RECT 110.230 173.120 110.510 173.400 ;
        RECT 112.205 173.175 112.485 173.455 ;
        RECT 112.605 173.175 112.885 173.455 ;
        RECT 88.640 172.665 88.920 172.945 ;
        RECT 108.355 172.745 108.635 173.025 ;
        RECT 108.755 172.745 109.035 173.025 ;
        RECT 110.230 172.720 110.510 173.000 ;
        RECT 112.205 172.745 112.485 173.025 ;
        RECT 112.605 172.745 112.885 173.025 ;
        RECT 108.355 172.315 108.635 172.595 ;
        RECT 108.755 172.315 109.035 172.595 ;
        RECT 112.205 172.315 112.485 172.595 ;
        RECT 112.605 172.315 112.885 172.595 ;
        RECT 108.355 171.455 108.635 171.735 ;
        RECT 108.755 171.455 109.035 171.735 ;
        RECT 112.205 171.455 112.485 171.735 ;
        RECT 112.605 171.455 112.885 171.735 ;
        RECT 108.355 170.595 108.635 170.875 ;
        RECT 108.755 170.595 109.035 170.875 ;
        RECT 112.205 170.595 112.485 170.875 ;
        RECT 112.605 170.595 112.885 170.875 ;
        RECT 108.355 170.165 108.635 170.445 ;
        RECT 108.755 170.165 109.035 170.445 ;
        RECT 110.230 170.285 110.510 170.565 ;
        RECT 112.205 170.165 112.485 170.445 ;
        RECT 112.605 170.165 112.885 170.445 ;
        RECT 108.355 169.735 108.635 170.015 ;
        RECT 108.755 169.735 109.035 170.015 ;
        RECT 110.230 169.885 110.510 170.165 ;
        RECT 108.355 169.065 108.635 169.345 ;
        RECT 108.755 169.065 109.035 169.345 ;
        RECT 112.205 169.735 112.485 170.015 ;
        RECT 112.605 169.735 112.885 170.015 ;
        RECT 112.205 169.065 112.485 169.345 ;
        RECT 112.605 169.065 112.885 169.345 ;
        RECT 116.810 167.700 117.090 167.980 ;
        RECT 116.810 167.300 117.090 167.580 ;
        RECT 116.810 166.900 117.090 167.180 ;
        RECT 123.705 166.180 123.985 166.460 ;
        RECT 123.705 165.780 123.985 166.060 ;
        RECT 123.705 165.380 123.985 165.660 ;
        RECT 109.815 164.695 110.095 164.975 ;
        RECT 111.185 164.695 111.465 164.975 ;
        RECT 112.555 164.695 112.835 164.975 ;
        RECT 123.020 164.655 123.300 164.935 ;
        RECT 109.815 164.025 110.095 164.305 ;
        RECT 111.185 164.025 111.465 164.305 ;
        RECT 112.555 164.025 112.835 164.305 ;
        RECT 123.020 164.025 123.300 164.305 ;
        RECT 109.815 161.745 110.095 162.025 ;
        RECT 111.185 161.745 111.465 162.025 ;
        RECT 112.555 161.745 112.835 162.025 ;
        RECT 123.020 161.745 123.300 162.025 ;
        RECT 124.390 164.655 124.670 164.935 ;
        RECT 124.390 164.025 124.670 164.305 ;
        RECT 124.390 161.745 124.670 162.025 ;
        RECT 109.815 159.465 110.095 159.745 ;
        RECT 111.185 159.465 111.465 159.745 ;
        RECT 112.555 159.465 112.835 159.745 ;
        RECT 123.020 157.185 123.300 157.465 ;
        RECT 109.815 154.905 110.095 155.185 ;
        RECT 78.070 154.360 78.350 154.640 ;
        RECT 78.470 154.360 78.750 154.640 ;
        RECT 78.870 154.360 79.150 154.640 ;
        RECT 104.665 154.360 104.945 154.640 ;
        RECT 105.065 154.360 105.345 154.640 ;
        RECT 105.465 154.360 105.745 154.640 ;
        RECT 80.170 153.260 80.450 153.540 ;
        RECT 80.570 153.260 80.850 153.540 ;
        RECT 80.970 153.260 81.250 153.540 ;
        RECT 106.260 153.420 106.540 153.700 ;
        RECT 106.260 153.020 106.540 153.300 ;
        RECT 111.185 154.905 111.465 155.185 ;
        RECT 124.390 157.185 124.670 157.465 ;
        RECT 112.555 154.905 112.835 155.185 ;
        RECT 106.260 152.620 106.540 152.900 ;
        RECT 123.020 152.625 123.300 152.905 ;
        RECT 63.195 151.930 63.475 152.210 ;
        RECT 63.595 151.930 63.875 152.210 ;
        RECT 63.995 151.930 64.275 152.210 ;
        RECT 71.335 151.885 71.615 152.165 ;
        RECT 57.310 151.445 57.590 151.725 ;
        RECT 57.710 151.445 57.990 151.725 ;
        RECT 60.900 151.445 61.180 151.725 ;
        RECT 61.300 151.445 61.580 151.725 ;
        RECT 65.515 151.445 65.795 151.725 ;
        RECT 71.335 151.485 71.615 151.765 ;
        RECT 71.335 151.085 71.615 151.365 ;
        RECT 60.900 150.775 61.180 151.055 ;
        RECT 61.300 150.775 61.580 151.055 ;
        RECT 65.515 150.775 65.795 151.055 ;
        RECT 87.175 151.885 87.455 152.165 ;
        RECT 94.515 151.930 94.795 152.210 ;
        RECT 94.915 151.930 95.195 152.210 ;
        RECT 95.315 151.930 95.595 152.210 ;
        RECT 87.175 151.485 87.455 151.765 ;
        RECT 92.995 151.445 93.275 151.725 ;
        RECT 97.210 151.445 97.490 151.725 ;
        RECT 97.610 151.445 97.890 151.725 ;
        RECT 100.800 151.445 101.080 151.725 ;
        RECT 101.200 151.445 101.480 151.725 ;
        RECT 87.175 151.085 87.455 151.365 ;
        RECT 92.995 150.775 93.275 151.055 ;
        RECT 97.210 150.775 97.490 151.055 ;
        RECT 97.610 150.775 97.890 151.055 ;
        RECT 109.815 150.345 110.095 150.625 ;
        RECT 60.900 149.995 61.180 150.275 ;
        RECT 61.300 149.995 61.580 150.275 ;
        RECT 65.515 149.995 65.795 150.275 ;
        RECT 92.995 149.995 93.275 150.275 ;
        RECT 97.210 149.995 97.490 150.275 ;
        RECT 97.610 149.995 97.890 150.275 ;
        RECT 63.195 149.605 63.475 149.885 ;
        RECT 60.900 149.215 61.180 149.495 ;
        RECT 61.300 149.215 61.580 149.495 ;
        RECT 95.315 149.605 95.595 149.885 ;
        RECT 63.195 149.205 63.475 149.485 ;
        RECT 65.515 149.215 65.795 149.495 ;
        RECT 92.995 149.215 93.275 149.495 ;
        RECT 63.195 148.805 63.475 149.085 ;
        RECT 95.315 149.205 95.595 149.485 ;
        RECT 97.210 149.215 97.490 149.495 ;
        RECT 97.610 149.215 97.890 149.495 ;
        RECT 95.315 148.805 95.595 149.085 ;
        RECT 111.185 150.345 111.465 150.625 ;
        RECT 124.390 152.625 124.670 152.905 ;
        RECT 112.555 150.345 112.835 150.625 ;
        RECT 123.020 148.065 123.300 148.345 ;
        RECT 62.710 146.935 62.990 147.215 ;
        RECT 63.110 146.935 63.390 147.215 ;
        RECT 63.790 146.890 64.070 147.170 ;
        RECT 63.790 146.490 64.070 146.770 ;
        RECT 72.160 146.890 72.440 147.170 ;
        RECT 63.790 146.090 64.070 146.370 ;
        RECT 72.160 146.490 72.440 146.770 ;
        RECT 72.160 146.090 72.440 146.370 ;
        RECT 86.350 146.890 86.630 147.170 ;
        RECT 86.350 146.490 86.630 146.770 ;
        RECT 94.720 146.890 95.000 147.170 ;
        RECT 95.400 146.935 95.680 147.215 ;
        RECT 95.800 146.935 96.080 147.215 ;
        RECT 86.350 146.090 86.630 146.370 ;
        RECT 94.720 146.490 95.000 146.770 ;
        RECT 94.720 146.090 95.000 146.370 ;
        RECT 109.815 145.785 110.095 146.065 ;
        RECT 60.900 144.655 61.180 144.935 ;
        RECT 61.300 144.655 61.580 144.935 ;
        RECT 65.515 144.655 65.795 144.935 ;
        RECT 92.995 144.655 93.275 144.935 ;
        RECT 97.210 144.655 97.490 144.935 ;
        RECT 97.610 144.655 97.890 144.935 ;
        RECT 60.900 143.875 61.180 144.155 ;
        RECT 61.300 143.875 61.580 144.155 ;
        RECT 65.515 143.875 65.795 144.155 ;
        RECT 92.995 143.875 93.275 144.155 ;
        RECT 97.210 143.875 97.490 144.155 ;
        RECT 97.610 143.875 97.890 144.155 ;
        RECT 111.185 145.785 111.465 146.065 ;
        RECT 124.390 148.065 124.670 148.345 ;
        RECT 112.555 145.785 112.835 146.065 ;
        RECT 123.020 143.505 123.300 143.785 ;
        RECT 60.900 143.095 61.180 143.375 ;
        RECT 61.300 143.095 61.580 143.375 ;
        RECT 65.515 143.095 65.795 143.375 ;
        RECT 92.995 143.095 93.275 143.375 ;
        RECT 97.210 143.095 97.490 143.375 ;
        RECT 97.610 143.095 97.890 143.375 ;
        RECT 73.670 142.725 73.950 143.005 ;
        RECT 76.410 142.725 76.690 143.005 ;
        RECT 82.100 142.725 82.380 143.005 ;
        RECT 84.840 142.725 85.120 143.005 ;
        RECT 60.900 142.315 61.180 142.595 ;
        RECT 61.300 142.315 61.580 142.595 ;
        RECT 65.515 142.425 65.795 142.705 ;
        RECT 92.995 142.425 93.275 142.705 ;
        RECT 73.670 142.095 73.950 142.375 ;
        RECT 57.310 141.535 57.590 141.815 ;
        RECT 57.710 141.535 57.990 141.815 ;
        RECT 76.410 141.695 76.690 141.975 ;
        RECT 78.205 141.865 78.485 142.145 ;
        RECT 57.310 139.255 57.590 139.535 ;
        RECT 57.710 139.255 57.990 139.535 ;
        RECT 78.205 141.465 78.485 141.745 ;
        RECT 78.205 141.065 78.485 141.345 ;
        RECT 80.305 141.865 80.585 142.145 ;
        RECT 84.840 142.095 85.120 142.375 ;
        RECT 97.210 142.315 97.490 142.595 ;
        RECT 97.610 142.315 97.890 142.595 ;
        RECT 80.305 141.465 80.585 141.745 ;
        RECT 82.100 141.695 82.380 141.975 ;
        RECT 100.800 141.535 101.080 141.815 ;
        RECT 101.200 141.535 101.480 141.815 ;
        RECT 80.305 141.065 80.585 141.345 ;
        RECT 75.080 139.735 75.360 140.015 ;
        RECT 62.710 139.255 62.990 139.535 ;
        RECT 63.110 139.255 63.390 139.535 ;
        RECT 75.080 139.335 75.360 139.615 ;
        RECT 83.430 139.735 83.710 140.015 ;
        RECT 83.430 139.335 83.710 139.615 ;
        RECT 95.400 139.255 95.680 139.535 ;
        RECT 95.800 139.255 96.080 139.535 ;
        RECT 65.515 138.235 65.795 138.515 ;
        RECT 69.320 138.235 69.600 138.515 ;
        RECT 69.720 138.235 70.000 138.515 ;
        RECT 76.410 138.415 76.690 138.695 ;
        RECT 82.100 138.415 82.380 138.695 ;
        RECT 88.790 138.235 89.070 138.515 ;
        RECT 89.190 138.235 89.470 138.515 ;
        RECT 92.995 138.235 93.275 138.515 ;
        RECT 65.515 137.565 65.795 137.845 ;
        RECT 69.320 137.565 69.600 137.845 ;
        RECT 69.720 137.565 70.000 137.845 ;
        RECT 88.790 137.565 89.070 137.845 ;
        RECT 89.190 137.565 89.470 137.845 ;
        RECT 92.995 137.565 93.275 137.845 ;
        RECT 57.310 136.975 57.590 137.255 ;
        RECT 57.710 136.975 57.990 137.255 ;
        RECT 72.160 137.210 72.440 137.490 ;
        RECT 57.310 134.695 57.590 134.975 ;
        RECT 57.710 134.695 57.990 134.975 ;
        RECT 72.160 136.810 72.440 137.090 ;
        RECT 65.515 136.285 65.795 136.565 ;
        RECT 69.320 136.285 69.600 136.565 ;
        RECT 69.720 136.285 70.000 136.565 ;
        RECT 72.160 136.410 72.440 136.690 ;
        RECT 65.515 135.005 65.795 135.285 ;
        RECT 69.320 135.005 69.600 135.285 ;
        RECT 69.720 135.005 70.000 135.285 ;
        RECT 62.710 134.695 62.990 134.975 ;
        RECT 63.110 134.695 63.390 134.975 ;
        RECT 67.705 134.205 67.985 134.485 ;
        RECT 67.705 133.805 67.985 134.085 ;
        RECT 67.705 133.405 67.985 133.685 ;
        RECT 86.350 137.210 86.630 137.490 ;
        RECT 109.815 141.225 110.095 141.505 ;
        RECT 100.800 139.255 101.080 139.535 ;
        RECT 101.200 139.255 101.480 139.535 ;
        RECT 111.185 141.225 111.465 141.505 ;
        RECT 124.390 143.505 124.670 143.785 ;
        RECT 112.555 141.225 112.835 141.505 ;
        RECT 123.020 138.945 123.300 139.225 ;
        RECT 86.350 136.810 86.630 137.090 ;
        RECT 100.800 136.975 101.080 137.255 ;
        RECT 101.200 136.975 101.480 137.255 ;
        RECT 86.350 136.410 86.630 136.690 ;
        RECT 75.080 135.175 75.360 135.455 ;
        RECT 76.410 135.135 76.690 135.415 ;
        RECT 82.100 135.135 82.380 135.415 ;
        RECT 83.430 135.175 83.710 135.455 ;
        RECT 75.080 134.775 75.360 135.055 ;
        RECT 83.430 134.775 83.710 135.055 ;
        RECT 88.790 136.285 89.070 136.565 ;
        RECT 89.190 136.285 89.470 136.565 ;
        RECT 92.995 136.285 93.275 136.565 ;
        RECT 88.790 135.005 89.070 135.285 ;
        RECT 89.190 135.005 89.470 135.285 ;
        RECT 92.995 135.005 93.275 135.285 ;
        RECT 90.805 134.205 91.085 134.485 ;
        RECT 90.805 133.805 91.085 134.085 ;
        RECT 95.400 134.695 95.680 134.975 ;
        RECT 95.800 134.695 96.080 134.975 ;
        RECT 90.805 133.405 91.085 133.685 ;
        RECT 124.390 138.945 124.670 139.225 ;
        RECT 109.815 136.665 110.095 136.945 ;
        RECT 111.185 136.665 111.465 136.945 ;
        RECT 112.555 136.665 112.835 136.945 ;
        RECT 100.800 134.695 101.080 134.975 ;
        RECT 101.200 134.695 101.480 134.975 ;
        RECT 123.020 134.385 123.300 134.665 ;
        RECT 57.310 132.415 57.590 132.695 ;
        RECT 57.710 132.415 57.990 132.695 ;
        RECT 100.800 132.415 101.080 132.695 ;
        RECT 101.200 132.415 101.480 132.695 ;
        RECT 57.310 130.135 57.590 130.415 ;
        RECT 57.710 130.135 57.990 130.415 ;
        RECT 56.125 128.675 56.405 128.955 ;
        RECT 56.125 128.275 56.405 128.555 ;
        RECT 56.125 127.875 56.405 128.155 ;
        RECT 67.025 132.045 67.305 132.325 ;
        RECT 67.025 131.645 67.305 131.925 ;
        RECT 91.485 132.045 91.765 132.325 ;
        RECT 67.025 131.245 67.305 131.525 ;
        RECT 91.485 131.645 91.765 131.925 ;
        RECT 91.485 131.245 91.765 131.525 ;
        RECT 65.515 130.445 65.795 130.725 ;
        RECT 69.320 130.445 69.600 130.725 ;
        RECT 69.720 130.445 70.000 130.725 ;
        RECT 75.080 130.615 75.360 130.895 ;
        RECT 62.710 130.135 62.990 130.415 ;
        RECT 63.110 130.135 63.390 130.415 ;
        RECT 75.080 130.215 75.360 130.495 ;
        RECT 83.430 130.615 83.710 130.895 ;
        RECT 83.430 130.215 83.710 130.495 ;
        RECT 88.790 130.445 89.070 130.725 ;
        RECT 89.190 130.445 89.470 130.725 ;
        RECT 92.995 130.445 93.275 130.725 ;
        RECT 95.400 130.135 95.680 130.415 ;
        RECT 95.800 130.135 96.080 130.415 ;
        RECT 65.515 129.165 65.795 129.445 ;
        RECT 69.320 129.165 69.600 129.445 ;
        RECT 69.720 129.165 70.000 129.445 ;
        RECT 73.670 129.135 73.950 129.415 ;
        RECT 84.840 129.135 85.120 129.415 ;
        RECT 88.790 129.165 89.070 129.445 ;
        RECT 89.190 129.165 89.470 129.445 ;
        RECT 92.995 129.165 93.275 129.445 ;
        RECT 75.080 128.255 75.360 128.535 ;
        RECT 65.515 127.885 65.795 128.165 ;
        RECT 69.320 127.885 69.600 128.165 ;
        RECT 69.720 127.885 70.000 128.165 ;
        RECT 83.430 128.255 83.710 128.535 ;
        RECT 73.670 127.855 73.950 128.135 ;
        RECT 75.080 127.855 75.360 128.135 ;
        RECT 83.430 127.855 83.710 128.135 ;
        RECT 84.840 127.855 85.120 128.135 ;
        RECT 88.790 127.885 89.070 128.165 ;
        RECT 89.190 127.885 89.470 128.165 ;
        RECT 92.995 127.885 93.275 128.165 ;
        RECT 109.815 132.105 110.095 132.385 ;
        RECT 111.185 132.105 111.465 132.385 ;
        RECT 112.555 132.105 112.835 132.385 ;
        RECT 100.800 130.135 101.080 130.415 ;
        RECT 101.200 130.135 101.480 130.415 ;
        RECT 124.390 134.385 124.670 134.665 ;
        RECT 123.020 129.825 123.300 130.105 ;
        RECT 102.385 128.675 102.665 128.955 ;
        RECT 102.385 128.275 102.665 128.555 ;
        RECT 102.385 127.875 102.665 128.155 ;
        RECT 57.310 125.575 57.590 125.855 ;
        RECT 57.710 125.575 57.990 125.855 ;
        RECT 75.080 127.455 75.360 127.735 ;
        RECT 83.430 127.455 83.710 127.735 ;
        RECT 65.515 126.605 65.795 126.885 ;
        RECT 69.320 126.605 69.600 126.885 ;
        RECT 69.720 126.605 70.000 126.885 ;
        RECT 73.670 126.575 73.950 126.855 ;
        RECT 77.510 126.495 77.790 126.775 ;
        RECT 77.510 126.095 77.790 126.375 ;
        RECT 81.000 126.495 81.280 126.775 ;
        RECT 84.840 126.575 85.120 126.855 ;
        RECT 88.790 126.605 89.070 126.885 ;
        RECT 89.190 126.605 89.470 126.885 ;
        RECT 92.995 126.605 93.275 126.885 ;
        RECT 81.000 126.095 81.280 126.375 ;
        RECT 62.710 125.575 62.990 125.855 ;
        RECT 63.110 125.575 63.390 125.855 ;
        RECT 65.515 125.325 65.795 125.605 ;
        RECT 69.320 125.325 69.600 125.605 ;
        RECT 69.720 125.325 70.000 125.605 ;
        RECT 75.080 125.495 75.360 125.775 ;
        RECT 75.080 125.095 75.360 125.375 ;
        RECT 83.430 125.495 83.710 125.775 ;
        RECT 83.430 125.095 83.710 125.375 ;
        RECT 88.790 125.325 89.070 125.605 ;
        RECT 89.190 125.325 89.470 125.605 ;
        RECT 92.995 125.325 93.275 125.605 ;
        RECT 95.400 125.575 95.680 125.855 ;
        RECT 95.800 125.575 96.080 125.855 ;
        RECT 63.790 123.890 64.070 124.170 ;
        RECT 57.310 123.295 57.590 123.575 ;
        RECT 57.710 123.295 57.990 123.575 ;
        RECT 63.110 123.445 63.390 123.725 ;
        RECT 63.790 123.490 64.070 123.770 ;
        RECT 94.720 123.890 95.000 124.170 ;
        RECT 57.310 121.015 57.590 121.295 ;
        RECT 57.710 121.015 57.990 121.295 ;
        RECT 63.110 123.045 63.390 123.325 ;
        RECT 63.790 123.090 64.070 123.370 ;
        RECT 94.720 123.490 95.000 123.770 ;
        RECT 63.110 122.645 63.390 122.925 ;
        RECT 71.335 122.890 71.615 123.170 ;
        RECT 71.335 122.490 71.615 122.770 ;
        RECT 71.335 122.090 71.615 122.370 ;
        RECT 71.335 121.690 71.615 121.970 ;
        RECT 62.710 121.015 62.990 121.295 ;
        RECT 63.110 121.015 63.390 121.295 ;
        RECT 65.515 120.765 65.795 121.045 ;
        RECT 69.320 120.765 69.600 121.045 ;
        RECT 69.720 120.765 70.000 121.045 ;
        RECT 65.515 119.485 65.795 119.765 ;
        RECT 69.320 119.485 69.600 119.765 ;
        RECT 69.720 119.485 70.000 119.765 ;
        RECT 57.310 118.735 57.590 119.015 ;
        RECT 57.710 118.735 57.990 119.015 ;
        RECT 87.175 122.890 87.455 123.170 ;
        RECT 94.720 123.090 95.000 123.370 ;
        RECT 95.400 123.445 95.680 123.725 ;
        RECT 109.815 127.545 110.095 127.825 ;
        RECT 111.185 127.545 111.465 127.825 ;
        RECT 112.555 127.545 112.835 127.825 ;
        RECT 100.800 125.575 101.080 125.855 ;
        RECT 101.200 125.575 101.480 125.855 ;
        RECT 124.390 129.825 124.670 130.105 ;
        RECT 123.020 125.265 123.300 125.545 ;
        RECT 124.390 125.265 124.670 125.545 ;
        RECT 95.400 123.045 95.680 123.325 ;
        RECT 100.800 123.295 101.080 123.575 ;
        RECT 101.200 123.295 101.480 123.575 ;
        RECT 87.175 122.490 87.455 122.770 ;
        RECT 95.400 122.645 95.680 122.925 ;
        RECT 87.175 122.090 87.455 122.370 ;
        RECT 87.175 121.690 87.455 121.970 ;
        RECT 75.080 120.935 75.360 121.215 ;
        RECT 83.430 120.935 83.710 121.215 ;
        RECT 75.080 120.535 75.360 120.815 ;
        RECT 76.410 120.575 76.690 120.855 ;
        RECT 82.100 120.575 82.380 120.855 ;
        RECT 83.430 120.535 83.710 120.815 ;
        RECT 88.790 120.765 89.070 121.045 ;
        RECT 89.190 120.765 89.470 121.045 ;
        RECT 92.995 120.765 93.275 121.045 ;
        RECT 95.400 121.015 95.680 121.295 ;
        RECT 95.800 121.015 96.080 121.295 ;
        RECT 88.790 119.485 89.070 119.765 ;
        RECT 89.190 119.485 89.470 119.765 ;
        RECT 92.995 119.485 93.275 119.765 ;
        RECT 109.815 122.985 110.095 123.265 ;
        RECT 111.185 122.985 111.465 123.265 ;
        RECT 112.555 122.985 112.835 123.265 ;
        RECT 100.800 121.015 101.080 121.295 ;
        RECT 101.200 121.015 101.480 121.295 ;
        RECT 100.800 118.735 101.080 119.015 ;
        RECT 101.200 118.735 101.480 119.015 ;
        RECT 57.310 116.455 57.590 116.735 ;
        RECT 57.710 116.455 57.990 116.735 ;
        RECT 65.515 118.205 65.795 118.485 ;
        RECT 69.320 118.205 69.600 118.485 ;
        RECT 69.720 118.205 70.000 118.485 ;
        RECT 88.790 118.205 89.070 118.485 ;
        RECT 89.190 118.205 89.470 118.485 ;
        RECT 92.995 118.205 93.275 118.485 ;
        RECT 65.515 117.535 65.795 117.815 ;
        RECT 69.320 117.535 69.600 117.815 ;
        RECT 69.720 117.535 70.000 117.815 ;
        RECT 76.410 117.295 76.690 117.575 ;
        RECT 82.100 117.295 82.380 117.575 ;
        RECT 88.790 117.535 89.070 117.815 ;
        RECT 89.190 117.535 89.470 117.815 ;
        RECT 92.995 117.535 93.275 117.815 ;
        RECT 62.710 116.455 62.990 116.735 ;
        RECT 63.110 116.455 63.390 116.735 ;
        RECT 75.080 116.375 75.360 116.655 ;
        RECT 75.080 115.975 75.360 116.255 ;
        RECT 83.430 116.375 83.710 116.655 ;
        RECT 95.400 116.455 95.680 116.735 ;
        RECT 95.800 116.455 96.080 116.735 ;
        RECT 83.430 115.975 83.710 116.255 ;
        RECT 78.925 114.645 79.205 114.925 ;
        RECT 79.325 114.645 79.605 114.925 ;
        RECT 79.725 114.645 80.005 114.925 ;
        RECT 109.815 118.425 110.095 118.705 ;
        RECT 111.185 118.425 111.465 118.705 ;
        RECT 112.555 118.425 112.835 118.705 ;
        RECT 100.800 116.455 101.080 116.735 ;
        RECT 101.200 116.455 101.480 116.735 ;
        RECT 123.020 120.705 123.300 120.985 ;
        RECT 124.390 120.705 124.670 120.985 ;
        RECT 115.400 117.105 115.680 117.385 ;
        RECT 115.400 116.705 115.680 116.985 ;
        RECT 117.740 116.445 118.020 116.725 ;
        RECT 57.310 114.175 57.590 114.455 ;
        RECT 57.710 114.175 57.990 114.455 ;
        RECT 76.410 114.015 76.690 114.295 ;
        RECT 82.100 114.015 82.380 114.295 ;
        RECT 100.800 114.175 101.080 114.455 ;
        RECT 101.200 114.175 101.480 114.455 ;
        RECT 60.900 113.395 61.180 113.675 ;
        RECT 61.300 113.395 61.580 113.675 ;
        RECT 73.670 113.615 73.950 113.895 ;
        RECT 84.840 113.615 85.120 113.895 ;
        RECT 109.815 113.865 110.095 114.145 ;
        RECT 111.185 113.865 111.465 114.145 ;
        RECT 112.555 113.865 112.835 114.145 ;
        RECT 64.475 113.285 64.755 113.565 ;
        RECT 64.875 113.285 65.155 113.565 ;
        RECT 69.225 113.285 69.505 113.565 ;
        RECT 89.285 113.285 89.565 113.565 ;
        RECT 93.635 113.285 93.915 113.565 ;
        RECT 94.035 113.285 94.315 113.565 ;
        RECT 97.210 113.395 97.490 113.675 ;
        RECT 97.610 113.395 97.890 113.675 ;
        RECT 73.670 112.985 73.950 113.265 ;
        RECT 76.410 112.985 76.690 113.265 ;
        RECT 82.100 112.985 82.380 113.265 ;
        RECT 84.840 112.985 85.120 113.265 ;
        RECT 60.900 112.615 61.180 112.895 ;
        RECT 61.300 112.615 61.580 112.895 ;
        RECT 64.475 112.615 64.755 112.895 ;
        RECT 64.875 112.615 65.155 112.895 ;
        RECT 69.225 112.615 69.505 112.895 ;
        RECT 89.285 112.615 89.565 112.895 ;
        RECT 93.635 112.615 93.915 112.895 ;
        RECT 94.035 112.615 94.315 112.895 ;
        RECT 97.210 112.615 97.490 112.895 ;
        RECT 97.610 112.615 97.890 112.895 ;
        RECT 57.310 111.945 57.590 112.225 ;
        RECT 57.710 111.945 57.990 112.225 ;
        RECT 60.900 111.945 61.180 112.225 ;
        RECT 61.300 111.945 61.580 112.225 ;
        RECT 97.210 111.945 97.490 112.225 ;
        RECT 97.610 111.945 97.890 112.225 ;
        RECT 100.800 111.945 101.080 112.225 ;
        RECT 101.200 111.945 101.480 112.225 ;
        RECT 117.740 116.045 118.020 116.325 ;
        RECT 117.740 115.645 118.020 115.925 ;
        RECT 117.740 115.245 118.020 115.525 ;
        RECT 117.740 114.845 118.020 115.125 ;
        RECT 117.740 114.445 118.020 114.725 ;
        RECT 117.740 114.045 118.020 114.325 ;
        RECT 117.740 113.645 118.020 113.925 ;
        RECT 120.380 114.200 120.660 114.480 ;
        RECT 120.380 113.800 120.660 114.080 ;
        RECT 117.740 113.245 118.020 113.525 ;
        RECT 120.380 113.400 120.660 113.680 ;
        RECT 123.020 116.145 123.300 116.425 ;
        RECT 124.390 116.145 124.670 116.425 ;
        RECT 117.740 112.845 118.020 113.125 ;
        RECT 117.740 112.445 118.020 112.725 ;
        RECT 117.740 112.045 118.020 112.325 ;
        RECT 117.740 111.645 118.020 111.925 ;
        RECT 64.475 110.335 64.755 110.615 ;
        RECT 64.875 110.335 65.155 110.615 ;
        RECT 69.225 110.335 69.505 110.615 ;
        RECT 89.285 110.335 89.565 110.615 ;
        RECT 93.635 110.335 93.915 110.615 ;
        RECT 94.035 110.335 94.315 110.615 ;
        RECT 109.815 109.305 110.095 109.585 ;
        RECT 111.185 109.305 111.465 109.585 ;
        RECT 112.555 109.305 112.835 109.585 ;
        RECT 64.475 108.055 64.755 108.335 ;
        RECT 64.875 108.055 65.155 108.335 ;
        RECT 69.225 108.055 69.505 108.335 ;
        RECT 89.285 108.055 89.565 108.335 ;
        RECT 93.635 108.055 93.915 108.335 ;
        RECT 94.035 108.055 94.315 108.335 ;
        RECT 67.025 107.700 67.305 107.980 ;
        RECT 67.025 107.300 67.305 107.580 ;
        RECT 67.025 106.900 67.305 107.180 ;
        RECT 67.705 107.700 67.985 107.980 ;
        RECT 67.705 107.300 67.985 107.580 ;
        RECT 67.705 106.900 67.985 107.180 ;
        RECT 90.805 107.700 91.085 107.980 ;
        RECT 90.805 107.300 91.085 107.580 ;
        RECT 90.805 106.900 91.085 107.180 ;
        RECT 91.485 107.700 91.765 107.980 ;
        RECT 91.485 107.300 91.765 107.580 ;
        RECT 117.740 111.245 118.020 111.525 ;
        RECT 116.810 110.555 117.090 110.835 ;
        RECT 116.810 110.155 117.090 110.435 ;
        RECT 91.485 106.900 91.765 107.180 ;
        RECT 109.815 104.745 110.095 105.025 ;
        RECT 111.185 104.745 111.465 105.025 ;
        RECT 112.555 104.745 112.835 105.025 ;
        RECT 64.475 103.495 64.755 103.775 ;
        RECT 64.875 103.495 65.155 103.775 ;
        RECT 69.225 103.495 69.505 103.775 ;
        RECT 89.285 103.495 89.565 103.775 ;
        RECT 93.635 103.495 93.915 103.775 ;
        RECT 94.035 103.495 94.315 103.775 ;
        RECT 114.310 100.945 114.590 101.225 ;
        RECT 114.310 100.545 114.590 100.825 ;
        RECT 109.815 100.185 110.095 100.465 ;
        RECT 111.185 100.185 111.465 100.465 ;
        RECT 112.555 100.185 112.835 100.465 ;
        RECT 114.310 100.145 114.590 100.425 ;
        RECT 123.020 111.585 123.300 111.865 ;
        RECT 124.390 111.585 124.670 111.865 ;
        RECT 123.020 107.025 123.300 107.305 ;
        RECT 124.390 107.025 124.670 107.305 ;
        RECT 123.020 102.465 123.300 102.745 ;
        RECT 124.390 102.465 124.670 102.745 ;
        RECT 64.475 98.935 64.755 99.215 ;
        RECT 64.875 98.935 65.155 99.215 ;
        RECT 69.225 98.935 69.505 99.215 ;
        RECT 89.285 98.935 89.565 99.215 ;
        RECT 93.635 98.935 93.915 99.215 ;
        RECT 94.035 98.935 94.315 99.215 ;
        RECT 114.310 97.775 114.590 98.055 ;
        RECT 114.310 97.375 114.590 97.655 ;
        RECT 114.310 96.975 114.590 97.255 ;
        RECT 66.965 96.655 67.245 96.935 ;
        RECT 67.365 96.655 67.645 96.935 ;
        RECT 67.765 96.655 68.045 96.935 ;
        RECT 90.745 96.655 91.025 96.935 ;
        RECT 91.145 96.655 91.425 96.935 ;
        RECT 91.545 96.655 91.825 96.935 ;
        RECT 109.815 95.625 110.095 95.905 ;
        RECT 111.185 95.625 111.465 95.905 ;
        RECT 112.555 95.625 112.835 95.905 ;
        RECT 64.475 94.375 64.755 94.655 ;
        RECT 64.875 94.375 65.155 94.655 ;
        RECT 69.225 94.375 69.505 94.655 ;
        RECT 89.285 94.375 89.565 94.655 ;
        RECT 93.635 94.375 93.915 94.655 ;
        RECT 94.035 94.375 94.315 94.655 ;
        RECT 123.020 97.905 123.300 98.185 ;
        RECT 124.390 97.905 124.670 98.185 ;
        RECT 64.475 92.095 64.755 92.375 ;
        RECT 64.875 92.095 65.155 92.375 ;
        RECT 69.225 92.095 69.505 92.375 ;
        RECT 89.285 92.095 89.565 92.375 ;
        RECT 93.635 92.095 93.915 92.375 ;
        RECT 94.035 92.095 94.315 92.375 ;
        RECT 123.020 93.345 123.300 93.625 ;
        RECT 124.390 93.345 124.670 93.625 ;
        RECT 109.815 91.065 110.095 91.345 ;
        RECT 111.185 91.065 111.465 91.345 ;
        RECT 112.555 91.065 112.835 91.345 ;
        RECT 64.475 89.815 64.755 90.095 ;
        RECT 64.875 89.815 65.155 90.095 ;
        RECT 69.225 89.815 69.505 90.095 ;
        RECT 89.285 89.815 89.565 90.095 ;
        RECT 93.635 89.815 93.915 90.095 ;
        RECT 94.035 89.815 94.315 90.095 ;
        RECT 64.475 89.145 64.755 89.425 ;
        RECT 64.875 89.145 65.155 89.425 ;
        RECT 69.225 89.145 69.505 89.425 ;
        RECT 89.285 89.145 89.565 89.425 ;
        RECT 93.635 89.145 93.915 89.425 ;
        RECT 94.035 89.145 94.315 89.425 ;
        RECT 123.020 88.785 123.300 89.065 ;
        RECT 124.390 88.785 124.670 89.065 ;
        RECT 79.190 86.650 79.470 86.930 ;
        RECT 79.590 86.650 79.870 86.930 ;
        RECT 79.990 86.650 80.270 86.930 ;
        RECT 104.230 86.810 104.510 87.090 ;
        RECT 104.230 86.410 104.510 86.690 ;
        RECT 109.815 86.505 110.095 86.785 ;
        RECT 111.185 86.505 111.465 86.785 ;
        RECT 112.555 86.505 112.835 86.785 ;
        RECT 104.230 86.010 104.510 86.290 ;
        RECT 83.825 84.980 84.105 85.260 ;
        RECT 84.225 84.980 84.505 85.260 ;
        RECT 74.455 83.850 74.735 84.130 ;
        RECT 74.855 83.850 75.135 84.130 ;
        RECT 75.255 83.850 75.535 84.130 ;
        RECT 86.310 83.850 86.590 84.130 ;
        RECT 86.710 83.850 86.990 84.130 ;
        RECT 87.110 83.850 87.390 84.130 ;
        RECT 71.950 83.200 72.230 83.480 ;
        RECT 71.950 82.800 72.230 83.080 ;
        RECT 78.610 83.200 78.890 83.480 ;
        RECT 71.950 82.400 72.230 82.680 ;
        RECT 72.680 82.615 72.960 82.895 ;
        RECT 73.080 82.615 73.360 82.895 ;
        RECT 75.905 82.615 76.185 82.895 ;
        RECT 76.305 82.615 76.585 82.895 ;
        RECT 77.480 82.615 77.760 82.895 ;
        RECT 77.880 82.615 78.160 82.895 ;
        RECT 78.610 82.800 78.890 83.080 ;
        RECT 78.610 82.400 78.890 82.680 ;
        RECT 79.670 83.200 79.950 83.480 ;
        RECT 79.670 82.800 79.950 83.080 ;
        RECT 86.330 83.200 86.610 83.480 ;
        RECT 79.670 82.400 79.950 82.680 ;
        RECT 80.400 82.615 80.680 82.895 ;
        RECT 80.800 82.615 81.080 82.895 ;
        RECT 81.975 82.615 82.255 82.895 ;
        RECT 82.375 82.615 82.655 82.895 ;
        RECT 85.200 82.615 85.480 82.895 ;
        RECT 85.600 82.615 85.880 82.895 ;
        RECT 86.330 82.800 86.610 83.080 ;
        RECT 86.330 82.400 86.610 82.680 ;
        RECT 72.680 81.945 72.960 82.225 ;
        RECT 73.080 81.945 73.360 82.225 ;
        RECT 72.680 81.515 72.960 81.795 ;
        RECT 73.080 81.515 73.360 81.795 ;
        RECT 74.455 81.775 74.735 82.055 ;
        RECT 75.905 81.945 76.185 82.225 ;
        RECT 76.305 81.945 76.585 82.225 ;
        RECT 77.480 81.945 77.760 82.225 ;
        RECT 77.880 81.945 78.160 82.225 ;
        RECT 80.400 81.945 80.680 82.225 ;
        RECT 80.800 81.945 81.080 82.225 ;
        RECT 81.975 81.945 82.255 82.225 ;
        RECT 82.375 81.945 82.655 82.225 ;
        RECT 74.455 81.375 74.735 81.655 ;
        RECT 75.905 81.515 76.185 81.795 ;
        RECT 76.305 81.515 76.585 81.795 ;
        RECT 77.480 81.515 77.760 81.795 ;
        RECT 77.880 81.515 78.160 81.795 ;
        RECT 80.400 81.515 80.680 81.795 ;
        RECT 80.800 81.515 81.080 81.795 ;
        RECT 81.975 81.515 82.255 81.795 ;
        RECT 82.375 81.515 82.655 81.795 ;
        RECT 83.825 81.775 84.105 82.055 ;
        RECT 85.200 81.945 85.480 82.225 ;
        RECT 85.600 81.945 85.880 82.225 ;
        RECT 71.950 80.855 72.230 81.135 ;
        RECT 72.680 81.085 72.960 81.365 ;
        RECT 73.080 81.085 73.360 81.365 ;
        RECT 83.825 81.375 84.105 81.655 ;
        RECT 85.200 81.515 85.480 81.795 ;
        RECT 85.600 81.515 85.880 81.795 ;
        RECT 77.480 81.085 77.760 81.365 ;
        RECT 77.880 81.085 78.160 81.365 ;
        RECT 71.950 80.455 72.230 80.735 ;
        RECT 72.680 80.225 72.960 80.505 ;
        RECT 73.080 80.225 73.360 80.505 ;
        RECT 78.610 80.625 78.890 80.905 ;
        RECT 77.480 80.225 77.760 80.505 ;
        RECT 77.880 80.225 78.160 80.505 ;
        RECT 78.610 80.225 78.890 80.505 ;
        RECT 78.610 79.825 78.890 80.105 ;
        RECT 72.680 79.365 72.960 79.645 ;
        RECT 73.080 79.365 73.360 79.645 ;
        RECT 72.680 78.935 72.960 79.215 ;
        RECT 73.080 78.935 73.360 79.215 ;
        RECT 74.455 79.155 74.735 79.435 ;
        RECT 77.480 79.365 77.760 79.645 ;
        RECT 77.880 79.365 78.160 79.645 ;
        RECT 80.400 81.085 80.680 81.365 ;
        RECT 80.800 81.085 81.080 81.365 ;
        RECT 85.200 81.085 85.480 81.365 ;
        RECT 85.600 81.085 85.880 81.365 ;
        RECT 79.670 80.625 79.950 80.905 ;
        RECT 86.330 80.855 86.610 81.135 ;
        RECT 79.670 80.225 79.950 80.505 ;
        RECT 80.400 80.225 80.680 80.505 ;
        RECT 80.800 80.225 81.080 80.505 ;
        RECT 79.670 79.825 79.950 80.105 ;
        RECT 85.200 80.225 85.480 80.505 ;
        RECT 85.600 80.225 85.880 80.505 ;
        RECT 86.330 80.455 86.610 80.735 ;
        RECT 80.400 79.365 80.680 79.645 ;
        RECT 80.800 79.365 81.080 79.645 ;
        RECT 72.680 78.505 72.960 78.785 ;
        RECT 73.080 78.505 73.360 78.785 ;
        RECT 74.455 78.755 74.735 79.035 ;
        RECT 75.905 78.935 76.185 79.215 ;
        RECT 76.305 78.935 76.585 79.215 ;
        RECT 77.480 78.935 77.760 79.215 ;
        RECT 77.880 78.935 78.160 79.215 ;
        RECT 80.400 78.935 80.680 79.215 ;
        RECT 80.800 78.935 81.080 79.215 ;
        RECT 81.975 78.935 82.255 79.215 ;
        RECT 82.375 78.935 82.655 79.215 ;
        RECT 83.825 79.155 84.105 79.435 ;
        RECT 85.200 79.365 85.480 79.645 ;
        RECT 85.600 79.365 85.880 79.645 ;
        RECT 75.905 78.505 76.185 78.785 ;
        RECT 76.305 78.505 76.585 78.785 ;
        RECT 77.480 78.505 77.760 78.785 ;
        RECT 77.880 78.505 78.160 78.785 ;
        RECT 80.400 78.505 80.680 78.785 ;
        RECT 80.800 78.505 81.080 78.785 ;
        RECT 81.975 78.505 82.255 78.785 ;
        RECT 82.375 78.505 82.655 78.785 ;
        RECT 83.825 78.755 84.105 79.035 ;
        RECT 85.200 78.935 85.480 79.215 ;
        RECT 85.600 78.935 85.880 79.215 ;
        RECT 74.455 78.200 74.735 78.480 ;
        RECT 72.680 77.855 72.960 78.135 ;
        RECT 73.080 77.855 73.360 78.135 ;
        RECT 85.200 78.505 85.480 78.785 ;
        RECT 85.600 78.505 85.880 78.785 ;
        RECT 83.825 78.200 84.105 78.480 ;
        RECT 74.455 77.800 74.735 78.080 ;
        RECT 75.905 77.855 76.185 78.135 ;
        RECT 76.305 77.855 76.585 78.135 ;
        RECT 77.480 77.855 77.760 78.135 ;
        RECT 77.880 77.855 78.160 78.135 ;
        RECT 80.400 77.855 80.680 78.135 ;
        RECT 80.800 77.855 81.080 78.135 ;
        RECT 81.975 77.855 82.255 78.135 ;
        RECT 82.375 77.855 82.655 78.135 ;
        RECT 87.110 78.200 87.390 78.480 ;
        RECT 83.825 77.800 84.105 78.080 ;
        RECT 85.200 77.855 85.480 78.135 ;
        RECT 85.600 77.855 85.880 78.135 ;
        RECT 87.110 77.800 87.390 78.080 ;
        RECT 74.455 77.400 74.735 77.680 ;
        RECT 78.870 77.380 79.150 77.660 ;
        RECT 79.270 77.380 79.550 77.660 ;
        RECT 79.670 77.380 79.950 77.660 ;
        RECT 83.825 77.400 84.105 77.680 ;
        RECT 87.110 77.400 87.390 77.680 ;
        RECT 123.020 86.505 123.300 86.785 ;
        RECT 124.390 86.505 124.670 86.785 ;
        RECT 123.020 84.225 123.300 84.505 ;
        RECT 124.390 84.225 124.670 84.505 ;
        RECT 89.270 82.965 89.550 83.245 ;
        RECT 89.670 82.965 89.950 83.245 ;
        RECT 93.120 82.965 93.400 83.245 ;
        RECT 93.520 82.965 93.800 83.245 ;
        RECT 89.270 82.295 89.550 82.575 ;
        RECT 89.670 82.295 89.950 82.575 ;
        RECT 91.145 82.240 91.425 82.520 ;
        RECT 93.120 82.295 93.400 82.575 ;
        RECT 93.520 82.295 93.800 82.575 ;
        RECT 89.270 81.865 89.550 82.145 ;
        RECT 89.670 81.865 89.950 82.145 ;
        RECT 115.400 82.905 115.680 83.185 ;
        RECT 115.400 82.505 115.680 82.785 ;
        RECT 91.145 81.840 91.425 82.120 ;
        RECT 93.120 81.865 93.400 82.145 ;
        RECT 93.520 81.865 93.800 82.145 ;
        RECT 109.815 81.945 110.095 82.225 ;
        RECT 111.185 81.945 111.465 82.225 ;
        RECT 112.555 81.945 112.835 82.225 ;
        RECT 117.740 82.245 118.020 82.525 ;
        RECT 89.270 81.435 89.550 81.715 ;
        RECT 89.670 81.435 89.950 81.715 ;
        RECT 93.120 81.435 93.400 81.715 ;
        RECT 93.520 81.435 93.800 81.715 ;
        RECT 89.270 80.575 89.550 80.855 ;
        RECT 89.670 80.575 89.950 80.855 ;
        RECT 93.120 80.575 93.400 80.855 ;
        RECT 93.520 80.575 93.800 80.855 ;
        RECT 89.270 79.715 89.550 79.995 ;
        RECT 89.670 79.715 89.950 79.995 ;
        RECT 93.120 79.715 93.400 79.995 ;
        RECT 93.520 79.715 93.800 79.995 ;
        RECT 117.740 81.845 118.020 82.125 ;
        RECT 89.270 79.285 89.550 79.565 ;
        RECT 89.670 79.285 89.950 79.565 ;
        RECT 91.145 79.405 91.425 79.685 ;
        RECT 93.120 79.285 93.400 79.565 ;
        RECT 93.520 79.285 93.800 79.565 ;
        RECT 89.270 78.855 89.550 79.135 ;
        RECT 89.670 78.855 89.950 79.135 ;
        RECT 91.145 79.005 91.425 79.285 ;
        RECT 89.270 78.185 89.550 78.465 ;
        RECT 89.670 78.185 89.950 78.465 ;
        RECT 93.120 78.855 93.400 79.135 ;
        RECT 93.520 78.855 93.800 79.135 ;
        RECT 93.120 78.185 93.400 78.465 ;
        RECT 93.520 78.185 93.800 78.465 ;
        RECT 109.815 77.385 110.095 77.665 ;
        RECT 111.185 77.385 111.465 77.665 ;
        RECT 112.555 77.385 112.835 77.665 ;
        RECT 117.740 81.445 118.020 81.725 ;
        RECT 117.740 81.045 118.020 81.325 ;
        RECT 121.180 81.900 121.460 82.180 ;
        RECT 124.390 81.945 124.670 82.225 ;
        RECT 121.180 81.500 121.460 81.780 ;
        RECT 121.180 81.100 121.460 81.380 ;
        RECT 117.740 80.645 118.020 80.925 ;
        RECT 117.740 80.245 118.020 80.525 ;
        RECT 117.740 79.845 118.020 80.125 ;
        RECT 117.740 79.445 118.020 79.725 ;
        RECT 120.380 80.000 120.660 80.280 ;
        RECT 120.380 79.600 120.660 79.880 ;
        RECT 123.020 79.665 123.300 79.945 ;
        RECT 124.390 79.665 124.670 79.945 ;
        RECT 117.740 79.045 118.020 79.325 ;
        RECT 120.380 79.200 120.660 79.480 ;
        RECT 117.740 78.645 118.020 78.925 ;
        RECT 117.740 78.245 118.020 78.525 ;
        RECT 117.740 77.845 118.020 78.125 ;
        RECT 117.740 77.445 118.020 77.725 ;
        RECT 123.020 77.385 123.300 77.665 ;
        RECT 124.390 77.385 124.670 77.665 ;
        RECT 76.385 76.170 76.665 76.450 ;
        RECT 76.385 75.770 76.665 76.050 ;
        RECT 91.145 75.100 91.425 75.380 ;
        RECT 94.670 75.120 94.950 75.400 ;
        RECT 95.070 75.120 95.350 75.400 ;
        RECT 95.470 75.120 95.750 75.400 ;
        RECT 117.740 77.045 118.020 77.325 ;
        RECT 123.020 76.755 123.300 77.035 ;
        RECT 124.390 76.755 124.670 77.035 ;
        RECT 116.810 76.355 117.090 76.635 ;
        RECT 116.810 75.955 117.090 76.235 ;
        RECT 115.955 75.350 116.235 75.630 ;
        RECT 91.145 74.700 91.425 74.980 ;
        RECT 91.145 74.300 91.425 74.580 ;
        RECT 109.815 72.825 110.095 73.105 ;
        RECT 111.185 72.825 111.465 73.105 ;
        RECT 112.555 72.825 112.835 73.105 ;
        RECT 65.490 72.305 65.770 72.585 ;
        RECT 65.890 72.305 66.170 72.585 ;
        RECT 69.340 72.305 69.620 72.585 ;
        RECT 69.740 72.305 70.020 72.585 ;
        RECT 74.510 72.305 74.790 72.585 ;
        RECT 74.910 72.305 75.190 72.585 ;
        RECT 78.360 72.305 78.640 72.585 ;
        RECT 78.760 72.305 79.040 72.585 ;
        RECT 81.450 72.305 81.730 72.585 ;
        RECT 81.850 72.305 82.130 72.585 ;
        RECT 85.300 72.305 85.580 72.585 ;
        RECT 85.700 72.305 85.980 72.585 ;
        RECT 89.270 72.305 89.550 72.585 ;
        RECT 89.670 72.305 89.950 72.585 ;
        RECT 93.120 72.305 93.400 72.585 ;
        RECT 93.520 72.305 93.800 72.585 ;
        RECT 65.490 71.635 65.770 71.915 ;
        RECT 65.890 71.635 66.170 71.915 ;
        RECT 67.365 71.580 67.645 71.860 ;
        RECT 69.340 71.635 69.620 71.915 ;
        RECT 69.740 71.635 70.020 71.915 ;
        RECT 74.510 71.635 74.790 71.915 ;
        RECT 74.910 71.635 75.190 71.915 ;
        RECT 65.490 71.205 65.770 71.485 ;
        RECT 65.890 71.205 66.170 71.485 ;
        RECT 76.385 71.580 76.665 71.860 ;
        RECT 78.360 71.635 78.640 71.915 ;
        RECT 78.760 71.635 79.040 71.915 ;
        RECT 81.450 71.635 81.730 71.915 ;
        RECT 81.850 71.635 82.130 71.915 ;
        RECT 67.365 71.180 67.645 71.460 ;
        RECT 69.340 71.205 69.620 71.485 ;
        RECT 69.740 71.205 70.020 71.485 ;
        RECT 74.510 71.205 74.790 71.485 ;
        RECT 74.910 71.205 75.190 71.485 ;
        RECT 83.825 71.580 84.105 71.860 ;
        RECT 85.300 71.635 85.580 71.915 ;
        RECT 85.700 71.635 85.980 71.915 ;
        RECT 89.270 71.635 89.550 71.915 ;
        RECT 89.670 71.635 89.950 71.915 ;
        RECT 76.385 71.180 76.665 71.460 ;
        RECT 78.360 71.205 78.640 71.485 ;
        RECT 78.760 71.205 79.040 71.485 ;
        RECT 81.450 71.205 81.730 71.485 ;
        RECT 81.850 71.205 82.130 71.485 ;
        RECT 91.145 71.580 91.425 71.860 ;
        RECT 93.120 71.635 93.400 71.915 ;
        RECT 93.520 71.635 93.800 71.915 ;
        RECT 83.825 71.180 84.105 71.460 ;
        RECT 85.300 71.205 85.580 71.485 ;
        RECT 85.700 71.205 85.980 71.485 ;
        RECT 89.270 71.205 89.550 71.485 ;
        RECT 89.670 71.205 89.950 71.485 ;
        RECT 91.145 71.180 91.425 71.460 ;
        RECT 93.120 71.205 93.400 71.485 ;
        RECT 93.520 71.205 93.800 71.485 ;
        RECT 65.490 70.775 65.770 71.055 ;
        RECT 65.890 70.775 66.170 71.055 ;
        RECT 69.340 70.775 69.620 71.055 ;
        RECT 69.740 70.775 70.020 71.055 ;
        RECT 74.510 70.775 74.790 71.055 ;
        RECT 74.910 70.775 75.190 71.055 ;
        RECT 78.360 70.775 78.640 71.055 ;
        RECT 78.760 70.775 79.040 71.055 ;
        RECT 81.450 70.775 81.730 71.055 ;
        RECT 81.850 70.775 82.130 71.055 ;
        RECT 85.300 70.775 85.580 71.055 ;
        RECT 85.700 70.775 85.980 71.055 ;
        RECT 89.270 70.775 89.550 71.055 ;
        RECT 89.670 70.775 89.950 71.055 ;
        RECT 93.120 70.775 93.400 71.055 ;
        RECT 93.520 70.775 93.800 71.055 ;
        RECT 123.985 71.205 124.265 71.485 ;
        RECT 115.955 70.575 116.235 70.855 ;
        RECT 65.490 69.915 65.770 70.195 ;
        RECT 65.890 69.915 66.170 70.195 ;
        RECT 69.340 69.915 69.620 70.195 ;
        RECT 69.740 69.915 70.020 70.195 ;
        RECT 74.510 69.915 74.790 70.195 ;
        RECT 74.910 69.915 75.190 70.195 ;
        RECT 78.360 69.915 78.640 70.195 ;
        RECT 78.760 69.915 79.040 70.195 ;
        RECT 81.450 69.915 81.730 70.195 ;
        RECT 81.850 69.915 82.130 70.195 ;
        RECT 85.300 69.915 85.580 70.195 ;
        RECT 85.700 69.915 85.980 70.195 ;
        RECT 89.270 69.915 89.550 70.195 ;
        RECT 89.670 69.915 89.950 70.195 ;
        RECT 119.650 70.295 119.930 70.575 ;
        RECT 93.120 69.915 93.400 70.195 ;
        RECT 93.520 69.915 93.800 70.195 ;
        RECT 115.955 69.905 116.235 70.185 ;
        RECT 119.650 69.625 119.930 69.905 ;
        RECT 65.490 69.055 65.770 69.335 ;
        RECT 65.890 69.055 66.170 69.335 ;
        RECT 69.340 69.055 69.620 69.335 ;
        RECT 69.740 69.055 70.020 69.335 ;
        RECT 74.510 69.055 74.790 69.335 ;
        RECT 74.910 69.055 75.190 69.335 ;
        RECT 78.360 69.055 78.640 69.335 ;
        RECT 78.760 69.055 79.040 69.335 ;
        RECT 81.450 69.055 81.730 69.335 ;
        RECT 81.850 69.055 82.130 69.335 ;
        RECT 85.300 69.055 85.580 69.335 ;
        RECT 85.700 69.055 85.980 69.335 ;
        RECT 89.270 69.055 89.550 69.335 ;
        RECT 89.670 69.055 89.950 69.335 ;
        RECT 93.120 69.055 93.400 69.335 ;
        RECT 93.520 69.055 93.800 69.335 ;
        RECT 119.650 69.195 119.930 69.475 ;
        RECT 123.985 70.805 124.265 71.085 ;
        RECT 123.985 70.405 124.265 70.685 ;
        RECT 125.635 70.255 125.915 70.535 ;
        RECT 123.070 69.600 123.350 69.880 ;
        RECT 125.635 69.625 125.915 69.905 ;
        RECT 123.070 69.200 123.350 69.480 ;
        RECT 121.200 68.765 121.480 69.045 ;
        RECT 121.600 68.765 121.880 69.045 ;
        RECT 125.635 69.195 125.915 69.475 ;
        RECT 125.635 68.765 125.915 69.045 ;
        RECT 65.490 68.195 65.770 68.475 ;
        RECT 65.890 68.195 66.170 68.475 ;
        RECT 69.340 68.195 69.620 68.475 ;
        RECT 69.740 68.195 70.020 68.475 ;
        RECT 74.510 68.195 74.790 68.475 ;
        RECT 74.910 68.195 75.190 68.475 ;
        RECT 78.360 68.195 78.640 68.475 ;
        RECT 78.760 68.195 79.040 68.475 ;
        RECT 81.450 68.195 81.730 68.475 ;
        RECT 81.850 68.195 82.130 68.475 ;
        RECT 85.300 68.195 85.580 68.475 ;
        RECT 85.700 68.195 85.980 68.475 ;
        RECT 89.270 68.195 89.550 68.475 ;
        RECT 89.670 68.195 89.950 68.475 ;
        RECT 93.120 68.195 93.400 68.475 ;
        RECT 93.520 68.195 93.800 68.475 ;
        RECT 109.815 68.265 110.095 68.545 ;
        RECT 111.185 68.265 111.465 68.545 ;
        RECT 112.555 68.265 112.835 68.545 ;
        RECT 125.635 68.335 125.915 68.615 ;
        RECT 121.200 67.905 121.480 68.185 ;
        RECT 121.600 67.905 121.880 68.185 ;
        RECT 65.490 67.335 65.770 67.615 ;
        RECT 65.890 67.335 66.170 67.615 ;
        RECT 69.340 67.335 69.620 67.615 ;
        RECT 69.740 67.335 70.020 67.615 ;
        RECT 74.510 67.335 74.790 67.615 ;
        RECT 74.910 67.335 75.190 67.615 ;
        RECT 78.360 67.335 78.640 67.615 ;
        RECT 78.760 67.335 79.040 67.615 ;
        RECT 81.450 67.335 81.730 67.615 ;
        RECT 81.850 67.335 82.130 67.615 ;
        RECT 85.300 67.335 85.580 67.615 ;
        RECT 85.700 67.335 85.980 67.615 ;
        RECT 89.270 67.335 89.550 67.615 ;
        RECT 89.670 67.335 89.950 67.615 ;
        RECT 115.955 67.625 116.235 67.905 ;
        RECT 93.120 67.335 93.400 67.615 ;
        RECT 93.520 67.335 93.800 67.615 ;
        RECT 125.635 67.905 125.915 68.185 ;
        RECT 125.635 67.475 125.915 67.755 ;
        RECT 121.200 67.045 121.480 67.325 ;
        RECT 121.600 67.045 121.880 67.325 ;
        RECT 65.490 66.475 65.770 66.755 ;
        RECT 65.890 66.475 66.170 66.755 ;
        RECT 69.340 66.475 69.620 66.755 ;
        RECT 69.740 66.475 70.020 66.755 ;
        RECT 74.510 66.475 74.790 66.755 ;
        RECT 74.910 66.475 75.190 66.755 ;
        RECT 78.360 66.475 78.640 66.755 ;
        RECT 78.760 66.475 79.040 66.755 ;
        RECT 81.450 66.475 81.730 66.755 ;
        RECT 81.850 66.475 82.130 66.755 ;
        RECT 85.300 66.475 85.580 66.755 ;
        RECT 85.700 66.475 85.980 66.755 ;
        RECT 89.270 66.475 89.550 66.755 ;
        RECT 89.670 66.475 89.950 66.755 ;
        RECT 93.120 66.475 93.400 66.755 ;
        RECT 93.520 66.475 93.800 66.755 ;
        RECT 65.490 65.615 65.770 65.895 ;
        RECT 65.890 65.615 66.170 65.895 ;
        RECT 69.340 65.615 69.620 65.895 ;
        RECT 69.740 65.615 70.020 65.895 ;
        RECT 74.510 65.615 74.790 65.895 ;
        RECT 74.910 65.615 75.190 65.895 ;
        RECT 78.360 65.615 78.640 65.895 ;
        RECT 78.760 65.615 79.040 65.895 ;
        RECT 81.450 65.615 81.730 65.895 ;
        RECT 81.850 65.615 82.130 65.895 ;
        RECT 85.300 65.615 85.580 65.895 ;
        RECT 85.700 65.615 85.980 65.895 ;
        RECT 89.270 65.615 89.550 65.895 ;
        RECT 89.670 65.615 89.950 65.895 ;
        RECT 109.815 65.985 110.095 66.265 ;
        RECT 111.185 65.985 111.465 66.265 ;
        RECT 112.555 65.985 112.835 66.265 ;
        RECT 93.120 65.615 93.400 65.895 ;
        RECT 93.520 65.615 93.800 65.895 ;
        RECT 119.650 66.615 119.930 66.895 ;
        RECT 119.650 66.185 119.930 66.465 ;
        RECT 65.490 64.755 65.770 65.035 ;
        RECT 65.890 64.755 66.170 65.035 ;
        RECT 69.340 64.755 69.620 65.035 ;
        RECT 69.740 64.755 70.020 65.035 ;
        RECT 74.510 64.755 74.790 65.035 ;
        RECT 74.910 64.755 75.190 65.035 ;
        RECT 65.490 64.325 65.770 64.605 ;
        RECT 65.890 64.325 66.170 64.605 ;
        RECT 67.365 64.445 67.645 64.725 ;
        RECT 78.360 64.755 78.640 65.035 ;
        RECT 78.760 64.755 79.040 65.035 ;
        RECT 81.450 64.755 81.730 65.035 ;
        RECT 81.850 64.755 82.130 65.035 ;
        RECT 69.340 64.325 69.620 64.605 ;
        RECT 69.740 64.325 70.020 64.605 ;
        RECT 74.510 64.325 74.790 64.605 ;
        RECT 74.910 64.325 75.190 64.605 ;
        RECT 76.385 64.445 76.665 64.725 ;
        RECT 85.300 64.755 85.580 65.035 ;
        RECT 85.700 64.755 85.980 65.035 ;
        RECT 89.270 64.755 89.550 65.035 ;
        RECT 89.670 64.755 89.950 65.035 ;
        RECT 78.360 64.325 78.640 64.605 ;
        RECT 78.760 64.325 79.040 64.605 ;
        RECT 81.450 64.325 81.730 64.605 ;
        RECT 81.850 64.325 82.130 64.605 ;
        RECT 83.825 64.445 84.105 64.725 ;
        RECT 93.120 64.755 93.400 65.035 ;
        RECT 93.520 64.755 93.800 65.035 ;
        RECT 85.300 64.325 85.580 64.605 ;
        RECT 85.700 64.325 85.980 64.605 ;
        RECT 89.270 64.325 89.550 64.605 ;
        RECT 89.670 64.325 89.950 64.605 ;
        RECT 91.145 64.445 91.425 64.725 ;
        RECT 93.120 64.325 93.400 64.605 ;
        RECT 93.520 64.325 93.800 64.605 ;
        RECT 65.490 63.895 65.770 64.175 ;
        RECT 65.890 63.895 66.170 64.175 ;
        RECT 67.365 64.045 67.645 64.325 ;
        RECT 69.340 63.895 69.620 64.175 ;
        RECT 69.740 63.895 70.020 64.175 ;
        RECT 74.510 63.895 74.790 64.175 ;
        RECT 74.910 63.895 75.190 64.175 ;
        RECT 76.385 64.045 76.665 64.325 ;
        RECT 78.360 63.895 78.640 64.175 ;
        RECT 78.760 63.895 79.040 64.175 ;
        RECT 81.450 63.895 81.730 64.175 ;
        RECT 81.850 63.895 82.130 64.175 ;
        RECT 83.825 64.045 84.105 64.325 ;
        RECT 85.300 63.895 85.580 64.175 ;
        RECT 85.700 63.895 85.980 64.175 ;
        RECT 89.270 63.895 89.550 64.175 ;
        RECT 89.670 63.895 89.950 64.175 ;
        RECT 91.145 64.045 91.425 64.325 ;
        RECT 93.120 63.895 93.400 64.175 ;
        RECT 93.520 63.895 93.800 64.175 ;
        RECT 109.815 63.705 110.095 63.985 ;
        RECT 111.185 63.705 111.465 63.985 ;
        RECT 112.555 63.705 112.835 63.985 ;
        RECT 125.635 67.045 125.915 67.325 ;
        RECT 125.635 66.615 125.915 66.895 ;
        RECT 125.635 66.185 125.915 66.465 ;
        RECT 127.420 65.710 127.700 65.990 ;
        RECT 125.635 65.325 125.915 65.605 ;
        RECT 127.420 65.310 127.700 65.590 ;
        RECT 127.420 64.910 127.700 65.190 ;
        RECT 119.650 64.375 119.930 64.655 ;
        RECT 120.465 64.230 120.745 64.510 ;
        RECT 119.650 63.945 119.930 64.225 ;
        RECT 120.465 63.830 120.745 64.110 ;
        RECT 121.200 63.515 121.480 63.795 ;
        RECT 121.600 63.515 121.880 63.795 ;
        RECT 65.490 63.225 65.770 63.505 ;
        RECT 65.890 63.225 66.170 63.505 ;
        RECT 69.340 63.225 69.620 63.505 ;
        RECT 69.740 63.225 70.020 63.505 ;
        RECT 74.510 63.225 74.790 63.505 ;
        RECT 74.910 63.225 75.190 63.505 ;
        RECT 78.360 63.225 78.640 63.505 ;
        RECT 78.760 63.225 79.040 63.505 ;
        RECT 81.450 63.225 81.730 63.505 ;
        RECT 81.850 63.225 82.130 63.505 ;
        RECT 85.300 63.225 85.580 63.505 ;
        RECT 85.700 63.225 85.980 63.505 ;
        RECT 89.270 63.225 89.550 63.505 ;
        RECT 89.670 63.225 89.950 63.505 ;
        RECT 93.120 63.225 93.400 63.505 ;
        RECT 93.520 63.225 93.800 63.505 ;
        RECT 109.815 63.035 110.095 63.315 ;
        RECT 111.185 63.035 111.465 63.315 ;
        RECT 112.555 63.035 112.835 63.315 ;
        RECT 115.955 63.065 116.235 63.345 ;
        RECT 121.200 62.655 121.480 62.935 ;
        RECT 121.600 62.655 121.880 62.935 ;
        RECT 121.180 61.795 121.460 62.075 ;
        RECT 121.580 61.795 121.860 62.075 ;
        RECT 119.650 61.365 119.930 61.645 ;
        RECT 123.985 61.450 124.265 61.730 ;
        RECT 115.955 60.785 116.235 61.065 ;
        RECT 119.650 60.935 119.930 61.215 ;
        RECT 123.985 61.050 124.265 61.330 ;
        RECT 115.955 60.115 116.235 60.395 ;
        RECT 119.650 60.305 119.930 60.585 ;
        RECT 120.465 59.425 120.745 59.705 ;
        RECT 120.865 59.425 121.145 59.705 ;
        RECT 122.670 59.425 122.950 59.705 ;
        RECT 123.070 59.425 123.350 59.705 ;
        RECT 125.635 64.465 125.915 64.745 ;
        RECT 125.635 64.035 125.915 64.315 ;
        RECT 125.635 63.605 125.915 63.885 ;
        RECT 125.635 63.175 125.915 63.455 ;
        RECT 125.635 62.745 125.915 63.025 ;
        RECT 125.635 62.315 125.915 62.595 ;
        RECT 125.635 61.885 125.915 62.165 ;
        RECT 125.635 61.455 125.915 61.735 ;
        RECT 125.635 61.025 125.915 61.305 ;
        RECT 125.635 60.395 125.915 60.675 ;
        RECT 124.800 57.200 125.080 57.480 ;
        RECT 124.800 56.800 125.080 57.080 ;
        RECT 124.800 56.400 125.080 56.680 ;
        RECT 124.800 56.000 125.080 56.280 ;
        RECT 124.800 55.600 125.080 55.880 ;
        RECT 124.665 38.865 124.945 39.145 ;
        RECT 125.065 38.865 125.345 39.145 ;
        RECT 125.465 38.865 125.745 39.145 ;
        RECT 140.825 38.865 141.105 39.145 ;
        RECT 141.225 38.865 141.505 39.145 ;
        RECT 141.625 38.865 141.905 39.145 ;
        RECT 142.025 38.865 142.305 39.145 ;
        RECT 104.230 21.680 104.510 21.960 ;
        RECT 104.230 21.280 104.510 21.560 ;
        RECT 124.800 21.415 125.080 21.695 ;
        RECT 72.305 20.820 72.585 21.100 ;
        RECT 104.230 20.880 104.510 21.160 ;
        RECT 124.800 21.015 125.080 21.295 ;
        RECT 72.305 20.420 72.585 20.700 ;
        RECT 124.800 20.615 125.080 20.895 ;
        RECT 72.305 20.020 72.585 20.300 ;
        RECT 123.985 19.980 124.265 20.260 ;
        RECT 123.985 19.580 124.265 19.860 ;
        RECT 87.560 19.170 87.840 19.450 ;
        RECT 87.960 19.170 88.240 19.450 ;
        RECT 88.360 19.170 88.640 19.450 ;
        RECT 122.250 19.170 122.530 19.450 ;
        RECT 122.650 19.170 122.930 19.450 ;
        RECT 123.050 19.170 123.330 19.450 ;
        RECT 123.985 19.180 124.265 19.460 ;
        RECT 105.195 18.205 105.475 18.485 ;
        RECT 105.595 18.205 105.875 18.485 ;
        RECT 105.995 18.205 106.275 18.485 ;
        RECT 116.940 18.205 117.220 18.485 ;
        RECT 117.340 18.205 117.620 18.485 ;
        RECT 117.740 18.205 118.020 18.485 ;
        RECT 91.145 16.675 91.425 16.955 ;
        RECT 91.145 16.275 91.425 16.555 ;
        RECT 91.145 15.875 91.425 16.155 ;
        RECT 83.160 14.935 83.440 15.215 ;
        RECT 83.560 14.935 83.840 15.215 ;
        RECT 83.960 14.935 84.240 15.215 ;
        RECT 117.740 13.705 118.020 13.985 ;
        RECT 118.140 13.705 118.420 13.985 ;
        RECT 118.540 13.705 118.820 13.985 ;
        RECT 140.825 13.705 141.105 13.985 ;
        RECT 141.225 13.705 141.505 13.985 ;
        RECT 141.625 13.705 141.905 13.985 ;
        RECT 142.025 13.705 142.305 13.985 ;
        RECT 76.250 7.655 76.530 7.935 ;
        RECT 76.650 7.655 76.930 7.935 ;
        RECT 77.050 7.655 77.330 7.935 ;
        RECT 112.095 7.655 112.375 7.935 ;
        RECT 112.495 7.655 112.775 7.935 ;
        RECT 67.230 6.555 67.510 6.835 ;
        RECT 67.630 6.555 67.910 6.835 ;
        RECT 68.030 6.555 68.310 6.835 ;
        RECT 90.015 6.555 90.295 6.835 ;
        RECT 90.415 6.555 90.695 6.835 ;
        RECT 157.825 5.275 158.105 5.555 ;
        RECT 157.825 4.875 158.105 5.155 ;
        RECT 134.505 4.235 134.785 4.515 ;
        RECT 134.905 4.235 135.185 4.515 ;
        RECT 135.305 4.235 135.585 4.515 ;
        RECT 135.705 4.235 135.985 4.515 ;
        RECT 157.825 4.475 158.105 4.755 ;
        RECT 157.825 4.075 158.105 4.355 ;
      LAYER met3 ;
        RECT 3.980 219.260 81.585 220.760 ;
        RECT 127.395 211.800 128.525 212.130 ;
        RECT 142.980 211.800 144.160 212.130 ;
        RECT 115.375 210.970 116.505 211.300 ;
        RECT 106.100 206.445 107.230 207.045 ;
        RECT 84.910 173.720 85.290 174.870 ;
        RECT 88.590 172.620 88.970 173.770 ;
        RECT 1.000 168.955 55.500 171.955 ;
        RECT 49.000 64.410 52.000 163.435 ;
        RECT 52.500 59.680 55.500 168.955 ;
        RECT 78.045 154.200 79.175 154.800 ;
        RECT 63.170 151.905 64.300 152.235 ;
        RECT 56.100 127.830 56.430 139.435 ;
        RECT 57.150 89.435 58.150 151.850 ;
        RECT 60.740 111.820 61.740 151.850 ;
        RECT 63.170 148.760 63.500 151.905 ;
        RECT 62.685 146.910 63.415 147.240 ;
        RECT 63.085 139.560 63.415 146.910 ;
        RECT 62.685 139.230 63.415 139.560 ;
        RECT 63.085 135.000 63.415 139.230 ;
        RECT 62.685 134.670 63.415 135.000 ;
        RECT 63.085 130.440 63.415 134.670 ;
        RECT 62.685 130.110 63.415 130.440 ;
        RECT 62.685 125.550 63.415 125.880 ;
        RECT 63.085 121.320 63.415 125.550 ;
        RECT 63.765 123.045 64.095 147.215 ;
        RECT 62.685 120.990 63.415 121.320 ;
        RECT 63.085 116.760 63.415 120.990 ;
        RECT 62.685 116.430 63.415 116.760 ;
        RECT 65.405 114.435 65.905 151.850 ;
        RECT 64.315 89.020 65.315 113.635 ;
        RECT 67.000 106.875 67.330 134.535 ;
        RECT 67.680 106.875 68.010 134.530 ;
        RECT 69.160 117.410 70.160 138.640 ;
        RECT 66.940 96.630 68.070 96.960 ;
        RECT 67.340 84.100 67.670 96.630 ;
        RECT 69.115 89.020 69.615 115.435 ;
        RECT 71.310 112.225 71.640 152.210 ;
        RECT 72.135 136.385 72.465 147.215 ;
        RECT 73.560 91.435 74.060 143.075 ;
        RECT 75.055 115.950 75.385 140.040 ;
        RECT 72.595 89.435 74.060 91.435 ;
        RECT 76.300 89.435 76.800 143.075 ;
        RECT 78.045 141.040 78.645 154.200 ;
        RECT 80.145 153.700 80.745 154.800 ;
        RECT 104.640 154.200 105.770 154.800 ;
        RECT 80.145 153.100 81.275 153.700 ;
        RECT 80.145 141.040 80.745 153.100 ;
        RECT 77.460 125.875 77.840 126.995 ;
        RECT 80.950 125.875 81.330 126.995 ;
        RECT 78.900 114.620 80.030 114.950 ;
        RECT 67.340 83.770 72.255 84.100 ;
        RECT 65.330 63.160 66.330 72.710 ;
        RECT 67.340 71.145 67.670 83.770 ;
        RECT 71.925 80.430 72.255 83.770 ;
        RECT 1.000 56.680 55.500 59.680 ;
        RECT 67.205 6.995 67.805 64.815 ;
        RECT 69.180 63.160 70.180 79.435 ;
        RECT 72.595 77.830 73.445 89.435 ;
        RECT 79.165 87.090 79.765 114.620 ;
        RECT 81.990 89.435 82.490 143.075 ;
        RECT 83.405 115.950 83.735 140.040 ;
        RECT 84.730 91.435 85.230 143.075 ;
        RECT 86.325 136.385 86.655 147.215 ;
        RECT 87.150 112.225 87.480 152.210 ;
        RECT 94.490 151.905 95.620 152.235 ;
        RECT 88.630 117.410 89.630 138.640 ;
        RECT 84.730 89.435 85.965 91.435 ;
        RECT 79.165 86.490 80.295 87.090 ;
        RECT 83.800 84.955 84.530 85.285 ;
        RECT 74.430 83.825 75.560 84.155 ;
        RECT 74.430 81.285 74.760 83.825 ;
        RECT 74.430 77.355 74.760 79.575 ;
        RECT 75.820 77.830 76.670 82.920 ;
        RECT 77.395 77.830 78.245 82.920 ;
        RECT 78.585 79.640 78.915 83.525 ;
        RECT 79.645 77.685 79.975 83.550 ;
        RECT 80.315 79.435 81.165 82.920 ;
        RECT 81.890 79.435 82.740 82.920 ;
        RECT 83.800 81.285 84.130 84.955 ;
        RECT 80.315 77.830 82.740 79.435 ;
        RECT 78.845 77.355 79.975 77.685 ;
        RECT 76.360 75.090 76.690 76.540 ;
        RECT 72.280 74.760 76.690 75.090 ;
        RECT 72.280 19.975 72.610 74.760 ;
        RECT 74.350 63.160 75.350 72.710 ;
        RECT 76.360 71.145 76.690 74.760 ;
        RECT 76.225 8.095 76.825 64.815 ;
        RECT 78.200 63.160 79.200 72.710 ;
        RECT 81.290 63.160 82.290 77.830 ;
        RECT 83.800 75.090 84.130 79.575 ;
        RECT 85.115 77.830 85.965 89.435 ;
        RECT 89.175 89.020 89.675 115.435 ;
        RECT 90.780 106.875 91.110 134.530 ;
        RECT 91.460 106.875 91.790 134.535 ;
        RECT 92.885 114.435 93.385 151.850 ;
        RECT 95.290 148.760 95.620 151.905 ;
        RECT 94.695 123.045 95.025 147.215 ;
        RECT 95.375 146.910 96.105 147.240 ;
        RECT 95.375 139.560 95.705 146.910 ;
        RECT 95.375 139.230 96.105 139.560 ;
        RECT 95.375 135.000 95.705 139.230 ;
        RECT 95.375 134.670 96.105 135.000 ;
        RECT 95.375 130.440 95.705 134.670 ;
        RECT 95.375 130.110 96.105 130.440 ;
        RECT 95.375 125.550 96.105 125.880 ;
        RECT 95.375 121.320 95.705 125.550 ;
        RECT 95.375 120.990 96.105 121.320 ;
        RECT 95.375 116.760 95.705 120.990 ;
        RECT 95.375 116.430 96.105 116.760 ;
        RECT 90.720 96.630 91.850 96.960 ;
        RECT 91.120 84.460 91.450 96.630 ;
        RECT 93.475 89.020 94.475 113.635 ;
        RECT 97.050 111.820 98.050 151.850 ;
        RECT 100.640 89.435 101.640 151.850 ;
        RECT 102.360 127.830 102.690 139.435 ;
        RECT 86.285 83.825 87.415 84.155 ;
        RECT 86.305 80.430 86.635 83.525 ;
        RECT 87.085 77.355 87.415 83.825 ;
        RECT 91.120 84.130 95.775 84.460 ;
        RECT 83.800 74.760 87.845 75.090 ;
        RECT 83.800 71.145 84.130 74.760 ;
        RECT 83.665 15.375 84.265 64.815 ;
        RECT 85.140 63.160 86.140 72.710 ;
        RECT 87.515 19.475 87.845 74.760 ;
        RECT 89.110 63.160 90.110 83.370 ;
        RECT 91.120 81.805 91.450 84.130 ;
        RECT 91.120 78.325 91.450 79.775 ;
        RECT 91.120 71.145 91.450 75.425 ;
        RECT 87.515 19.145 88.665 19.475 ;
        RECT 90.985 15.850 91.585 64.815 ;
        RECT 92.960 63.160 93.960 83.370 ;
        RECT 95.445 75.425 95.775 84.130 ;
        RECT 94.645 75.095 95.775 75.425 ;
        RECT 104.070 20.855 104.670 87.115 ;
        RECT 105.170 18.645 105.770 154.200 ;
        RECT 106.100 19.150 106.700 206.445 ;
        RECT 115.375 175.950 115.705 210.970 ;
        RECT 120.355 210.140 121.485 210.470 ;
        RECT 117.715 207.940 118.845 208.540 ;
        RECT 110.195 175.620 115.705 175.950 ;
        RECT 108.195 169.000 109.195 174.250 ;
        RECT 110.195 173.985 110.525 175.620 ;
        RECT 110.195 173.655 110.535 173.985 ;
        RECT 110.205 172.685 110.535 173.655 ;
        RECT 110.205 169.205 110.535 170.655 ;
        RECT 112.045 169.000 113.045 174.250 ;
        RECT 108.195 167.380 108.895 169.000 ;
        RECT 107.250 166.680 108.895 167.380 ;
        RECT 107.250 161.435 107.950 166.680 ;
        RECT 109.605 63.010 110.305 165.000 ;
        RECT 110.975 63.010 111.675 165.000 ;
        RECT 112.345 63.010 113.045 169.000 ;
        RECT 114.285 96.845 114.615 101.280 ;
        RECT 115.375 76.305 115.705 175.620 ;
        RECT 116.785 75.920 117.115 207.045 ;
        RECT 117.715 111.080 118.045 207.940 ;
        RECT 115.745 60.090 116.445 75.655 ;
        RECT 117.715 18.645 118.045 82.690 ;
        RECT 120.355 79.175 120.685 210.140 ;
        RECT 123.680 209.040 124.410 209.640 ;
        RECT 123.680 165.255 124.010 209.040 ;
        RECT 119.440 65.570 120.140 70.600 ;
        RECT 121.155 69.070 121.485 82.225 ;
        RECT 122.810 76.730 123.510 164.960 ;
        RECT 124.180 73.925 124.880 164.960 ;
        RECT 124.180 73.225 126.125 73.925 ;
        RECT 121.155 68.740 121.905 69.070 ;
        RECT 121.155 68.210 121.485 68.740 ;
        RECT 121.155 67.880 121.905 68.210 ;
        RECT 121.155 67.350 121.485 67.880 ;
        RECT 121.155 67.020 121.905 67.350 ;
        RECT 119.440 60.280 120.140 65.230 ;
        RECT 120.440 59.730 120.770 64.715 ;
        RECT 121.155 63.820 121.485 67.020 ;
        RECT 121.155 63.490 121.905 63.820 ;
        RECT 121.155 62.960 121.485 63.490 ;
        RECT 121.155 62.630 121.905 62.960 ;
        RECT 121.155 62.100 121.485 62.630 ;
        RECT 121.155 61.770 121.885 62.100 ;
        RECT 123.045 59.730 123.375 70.055 ;
        RECT 120.440 59.400 121.170 59.730 ;
        RECT 122.645 59.400 123.375 59.730 ;
        RECT 123.045 19.475 123.375 59.400 ;
        RECT 122.225 19.145 123.375 19.475 ;
        RECT 105.170 18.045 106.300 18.645 ;
        RECT 116.915 18.045 118.045 18.645 ;
        RECT 123.045 18.045 123.375 19.145 ;
        RECT 123.960 18.045 124.290 71.530 ;
        RECT 125.425 60.370 126.125 73.225 ;
        RECT 124.640 39.305 125.240 57.560 ;
        RECT 124.640 38.705 125.770 39.305 ;
        RECT 124.640 18.045 125.240 38.705 ;
        RECT 127.395 18.045 127.725 211.800 ;
        RECT 146.655 210.140 147.835 210.470 ;
        RECT 140.605 207.940 142.530 208.540 ;
        RECT 129.470 184.540 153.530 207.140 ;
        RECT 129.470 159.245 153.530 181.845 ;
        RECT 129.470 135.445 153.530 158.045 ;
        RECT 129.470 111.645 153.530 134.245 ;
        RECT 129.470 87.845 153.530 110.445 ;
        RECT 129.470 64.045 153.530 86.645 ;
        RECT 129.470 40.245 153.530 62.845 ;
        RECT 140.605 38.705 142.530 39.305 ;
        RECT 83.135 14.775 84.265 15.375 ;
        RECT 117.715 14.145 118.045 18.045 ;
        RECT 129.470 14.945 153.530 37.545 ;
        RECT 117.715 13.545 118.845 14.145 ;
        RECT 140.605 13.545 142.530 14.145 ;
        RECT 76.225 7.495 77.355 8.095 ;
        RECT 111.875 7.495 113.000 8.095 ;
        RECT 67.205 6.395 68.335 6.995 ;
        RECT 89.795 6.395 90.920 6.995 ;
        RECT 134.480 4.075 136.010 4.675 ;
        RECT 90.320 1.810 90.920 3.750 ;
        RECT 112.400 1.810 113.000 3.750 ;
        RECT 134.480 1.810 135.080 3.750 ;
        RECT 156.565 1.810 157.165 209.665 ;
        RECT 157.665 4.050 158.265 211.325 ;
      LAYER via3 ;
        RECT 3.980 220.250 4.300 220.570 ;
        RECT 7.660 220.250 7.980 220.570 ;
        RECT 11.340 220.250 11.660 220.570 ;
        RECT 15.020 220.250 15.340 220.570 ;
        RECT 18.700 220.250 19.020 220.570 ;
        RECT 22.380 220.250 22.700 220.570 ;
        RECT 26.060 220.250 26.380 220.570 ;
        RECT 29.740 220.250 30.060 220.570 ;
        RECT 33.420 220.250 33.740 220.570 ;
        RECT 37.100 220.250 37.420 220.570 ;
        RECT 40.780 220.250 41.100 220.570 ;
        RECT 44.460 220.250 44.780 220.570 ;
        RECT 48.140 220.250 48.460 220.570 ;
        RECT 3.980 219.850 4.300 220.170 ;
        RECT 7.660 219.850 7.980 220.170 ;
        RECT 11.340 219.850 11.660 220.170 ;
        RECT 15.020 219.850 15.340 220.170 ;
        RECT 18.700 219.850 19.020 220.170 ;
        RECT 22.380 219.850 22.700 220.170 ;
        RECT 26.060 219.850 26.380 220.170 ;
        RECT 29.740 219.850 30.060 220.170 ;
        RECT 33.420 219.850 33.740 220.170 ;
        RECT 37.100 219.850 37.420 220.170 ;
        RECT 40.780 219.850 41.100 220.170 ;
        RECT 44.460 219.850 44.780 220.170 ;
        RECT 48.140 219.850 48.460 220.170 ;
        RECT 3.980 219.450 4.300 219.770 ;
        RECT 7.660 219.450 7.980 219.770 ;
        RECT 11.340 219.450 11.660 219.770 ;
        RECT 15.020 219.450 15.340 219.770 ;
        RECT 18.700 219.450 19.020 219.770 ;
        RECT 22.380 219.450 22.700 219.770 ;
        RECT 26.060 219.450 26.380 219.770 ;
        RECT 29.740 219.450 30.060 219.770 ;
        RECT 33.420 219.450 33.740 219.770 ;
        RECT 37.100 219.450 37.420 219.770 ;
        RECT 40.780 219.450 41.100 219.770 ;
        RECT 44.460 219.450 44.780 219.770 ;
        RECT 48.140 219.450 48.460 219.770 ;
        RECT 49.190 219.450 50.310 220.570 ;
        RECT 51.820 220.250 52.140 220.570 ;
        RECT 55.500 220.250 55.820 220.570 ;
        RECT 59.180 220.250 59.500 220.570 ;
        RECT 62.860 220.250 63.180 220.570 ;
        RECT 66.540 220.250 66.860 220.570 ;
        RECT 70.220 220.250 70.540 220.570 ;
        RECT 73.900 220.250 74.220 220.570 ;
        RECT 77.580 220.250 77.900 220.570 ;
        RECT 81.260 220.250 81.580 220.570 ;
        RECT 51.820 219.850 52.140 220.170 ;
        RECT 55.500 219.850 55.820 220.170 ;
        RECT 59.180 219.850 59.500 220.170 ;
        RECT 62.860 219.850 63.180 220.170 ;
        RECT 66.540 219.850 66.860 220.170 ;
        RECT 70.220 219.850 70.540 220.170 ;
        RECT 73.900 219.850 74.220 220.170 ;
        RECT 77.580 219.850 77.900 220.170 ;
        RECT 81.260 219.850 81.580 220.170 ;
        RECT 51.820 219.450 52.140 219.770 ;
        RECT 55.500 219.450 55.820 219.770 ;
        RECT 59.180 219.450 59.500 219.770 ;
        RECT 62.860 219.450 63.180 219.770 ;
        RECT 66.540 219.450 66.860 219.770 ;
        RECT 70.220 219.450 70.540 219.770 ;
        RECT 73.900 219.450 74.220 219.770 ;
        RECT 77.580 219.450 77.900 219.770 ;
        RECT 81.260 219.450 81.580 219.770 ;
        RECT 143.010 211.805 143.330 212.125 ;
        RECT 143.410 211.805 143.730 212.125 ;
        RECT 143.810 211.805 144.130 212.125 ;
        RECT 84.940 174.520 85.260 174.840 ;
        RECT 84.940 174.120 85.260 174.440 ;
        RECT 84.940 173.720 85.260 174.040 ;
        RECT 88.620 173.420 88.940 173.740 ;
        RECT 88.620 173.020 88.940 173.340 ;
        RECT 88.620 172.620 88.940 172.940 ;
        RECT 1.190 169.095 2.310 171.815 ;
        RECT 49.140 161.475 51.860 163.395 ;
        RECT 49.190 139.675 50.310 161.195 ;
        RECT 49.140 137.475 51.860 139.395 ;
        RECT 49.190 115.675 50.310 137.195 ;
        RECT 49.140 113.475 51.860 115.395 ;
        RECT 49.190 91.675 50.310 113.195 ;
        RECT 49.140 89.475 51.860 91.395 ;
        RECT 49.190 67.675 50.310 89.195 ;
        RECT 49.140 65.475 51.860 67.395 ;
        RECT 49.190 64.510 50.310 65.230 ;
        RECT 52.640 149.475 55.360 151.395 ;
        RECT 57.290 149.475 58.010 151.395 ;
        RECT 56.105 138.675 56.425 138.995 ;
        RECT 56.105 138.275 56.425 138.595 ;
        RECT 56.105 137.875 56.425 138.195 ;
        RECT 52.640 125.475 55.360 127.395 ;
        RECT 52.640 101.475 55.360 103.395 ;
        RECT 57.290 125.475 58.010 127.395 ;
        RECT 60.880 149.475 61.600 151.395 ;
        RECT 60.880 125.475 61.600 127.395 ;
        RECT 65.495 139.075 65.815 139.395 ;
        RECT 65.495 138.675 65.815 138.995 ;
        RECT 65.495 138.275 65.815 138.595 ;
        RECT 65.495 137.875 65.815 138.195 ;
        RECT 65.495 137.475 65.815 137.795 ;
        RECT 65.495 115.075 65.815 115.395 ;
        RECT 65.495 114.675 65.815 114.995 ;
        RECT 57.290 101.475 58.010 103.395 ;
        RECT 69.300 125.475 70.020 127.395 ;
        RECT 69.205 115.075 69.525 115.395 ;
        RECT 69.205 114.675 69.525 114.995 ;
        RECT 69.205 114.275 69.525 114.595 ;
        RECT 69.205 113.875 69.525 114.195 ;
        RECT 69.205 113.475 69.525 113.795 ;
        RECT 64.455 101.475 65.175 103.395 ;
        RECT 52.640 77.475 55.360 79.395 ;
        RECT 73.650 139.075 73.970 139.395 ;
        RECT 73.650 138.675 73.970 138.995 ;
        RECT 73.650 138.275 73.970 138.595 ;
        RECT 73.650 137.875 73.970 138.195 ;
        RECT 73.650 137.475 73.970 137.795 ;
        RECT 76.390 139.075 76.710 139.395 ;
        RECT 76.390 138.675 76.710 138.995 ;
        RECT 76.390 138.275 76.710 138.595 ;
        RECT 76.390 137.875 76.710 138.195 ;
        RECT 76.390 137.475 76.710 137.795 ;
        RECT 73.650 115.075 73.970 115.395 ;
        RECT 73.650 114.675 73.970 114.995 ;
        RECT 73.650 114.275 73.970 114.595 ;
        RECT 73.650 113.875 73.970 114.195 ;
        RECT 73.650 113.475 73.970 113.795 ;
        RECT 69.205 91.075 69.525 91.395 ;
        RECT 69.205 90.675 69.525 90.995 ;
        RECT 69.205 90.275 69.525 90.595 ;
        RECT 69.205 89.875 69.525 90.195 ;
        RECT 69.205 89.475 69.525 89.795 ;
        RECT 73.650 91.075 73.970 91.395 ;
        RECT 73.650 90.675 73.970 90.995 ;
        RECT 73.650 90.275 73.970 90.595 ;
        RECT 73.650 89.875 73.970 90.195 ;
        RECT 73.650 89.475 73.970 89.795 ;
        RECT 82.080 139.075 82.400 139.395 ;
        RECT 82.080 138.675 82.400 138.995 ;
        RECT 82.080 138.275 82.400 138.595 ;
        RECT 82.080 137.875 82.400 138.195 ;
        RECT 82.080 137.475 82.400 137.795 ;
        RECT 77.490 126.675 77.810 126.995 ;
        RECT 77.490 126.275 77.810 126.595 ;
        RECT 77.490 125.875 77.810 126.195 ;
        RECT 80.980 126.675 81.300 126.995 ;
        RECT 80.980 126.275 81.300 126.595 ;
        RECT 80.980 125.875 81.300 126.195 ;
        RECT 76.390 115.075 76.710 115.395 ;
        RECT 76.390 114.675 76.710 114.995 ;
        RECT 84.820 139.075 85.140 139.395 ;
        RECT 84.820 138.675 85.140 138.995 ;
        RECT 84.820 138.275 85.140 138.595 ;
        RECT 84.820 137.875 85.140 138.195 ;
        RECT 84.820 137.475 85.140 137.795 ;
        RECT 82.080 115.075 82.400 115.395 ;
        RECT 82.080 114.675 82.400 114.995 ;
        RECT 76.390 114.275 76.710 114.595 ;
        RECT 76.390 113.875 76.710 114.195 ;
        RECT 76.390 113.475 76.710 113.795 ;
        RECT 76.390 91.075 76.710 91.395 ;
        RECT 76.390 90.675 76.710 90.995 ;
        RECT 76.390 90.275 76.710 90.595 ;
        RECT 76.390 89.875 76.710 90.195 ;
        RECT 76.390 89.475 76.710 89.795 ;
        RECT 82.080 114.275 82.400 114.595 ;
        RECT 82.080 113.875 82.400 114.195 ;
        RECT 82.080 113.475 82.400 113.795 ;
        RECT 82.080 91.075 82.400 91.395 ;
        RECT 82.080 90.675 82.400 90.995 ;
        RECT 82.080 90.275 82.400 90.595 ;
        RECT 82.080 89.875 82.400 90.195 ;
        RECT 82.080 89.475 82.400 89.795 ;
        RECT 84.820 115.075 85.140 115.395 ;
        RECT 84.820 114.675 85.140 114.995 ;
        RECT 84.820 114.275 85.140 114.595 ;
        RECT 84.820 113.875 85.140 114.195 ;
        RECT 84.820 113.475 85.140 113.795 ;
        RECT 97.190 149.475 97.910 151.395 ;
        RECT 92.975 139.075 93.295 139.395 ;
        RECT 92.975 138.675 93.295 138.995 ;
        RECT 92.975 138.275 93.295 138.595 ;
        RECT 92.975 137.875 93.295 138.195 ;
        RECT 92.975 137.475 93.295 137.795 ;
        RECT 88.770 125.475 89.490 127.395 ;
        RECT 89.265 115.075 89.585 115.395 ;
        RECT 89.265 114.675 89.585 114.995 ;
        RECT 89.265 114.275 89.585 114.595 ;
        RECT 89.265 113.875 89.585 114.195 ;
        RECT 89.265 113.475 89.585 113.795 ;
        RECT 84.820 91.075 85.140 91.395 ;
        RECT 85.460 91.075 85.780 91.395 ;
        RECT 84.820 90.675 85.140 90.995 ;
        RECT 85.460 90.675 85.780 90.995 ;
        RECT 84.820 90.275 85.140 90.595 ;
        RECT 85.460 90.275 85.780 90.595 ;
        RECT 84.820 89.875 85.140 90.195 ;
        RECT 85.460 89.875 85.780 90.195 ;
        RECT 84.820 89.475 85.140 89.795 ;
        RECT 85.460 89.475 85.780 89.795 ;
        RECT 72.660 82.000 73.380 82.720 ;
        RECT 69.320 77.475 70.040 79.395 ;
        RECT 65.470 65.475 66.190 67.395 ;
        RECT 1.190 56.820 2.310 59.540 ;
        RECT 75.885 78.000 76.605 78.720 ;
        RECT 77.460 78.000 78.180 78.720 ;
        RECT 97.190 125.475 97.910 127.395 ;
        RECT 92.975 115.075 93.295 115.395 ;
        RECT 92.975 114.675 93.295 114.995 ;
        RECT 100.780 149.475 101.500 151.395 ;
        RECT 102.365 138.675 102.685 138.995 ;
        RECT 102.365 138.275 102.685 138.595 ;
        RECT 102.365 137.875 102.685 138.195 ;
        RECT 100.780 125.475 101.500 127.395 ;
        RECT 93.615 101.475 94.335 103.395 ;
        RECT 89.265 91.075 89.585 91.395 ;
        RECT 89.265 90.675 89.585 90.995 ;
        RECT 89.265 90.275 89.585 90.595 ;
        RECT 89.265 89.875 89.585 90.195 ;
        RECT 89.265 89.475 89.585 89.795 ;
        RECT 100.780 101.475 101.500 103.395 ;
        RECT 85.180 82.000 85.900 82.720 ;
        RECT 80.380 78.000 81.100 78.720 ;
        RECT 81.955 78.000 82.675 78.720 ;
        RECT 74.490 65.475 75.210 67.395 ;
        RECT 85.280 65.475 86.000 67.395 ;
        RECT 93.100 77.475 93.820 79.395 ;
        RECT 89.250 65.475 89.970 67.395 ;
        RECT 107.440 163.075 107.760 163.395 ;
        RECT 107.440 162.675 107.760 162.995 ;
        RECT 107.440 162.275 107.760 162.595 ;
        RECT 107.440 161.875 107.760 162.195 ;
        RECT 107.440 161.475 107.760 161.795 ;
        RECT 109.795 151.075 110.115 151.395 ;
        RECT 109.795 150.675 110.115 150.995 ;
        RECT 109.795 150.275 110.115 150.595 ;
        RECT 109.795 149.875 110.115 150.195 ;
        RECT 109.795 149.475 110.115 149.795 ;
        RECT 109.795 127.075 110.115 127.395 ;
        RECT 109.795 126.675 110.115 126.995 ;
        RECT 109.795 126.275 110.115 126.595 ;
        RECT 109.795 125.875 110.115 126.195 ;
        RECT 109.795 125.475 110.115 125.795 ;
        RECT 109.795 103.075 110.115 103.395 ;
        RECT 109.795 102.675 110.115 102.995 ;
        RECT 109.795 102.275 110.115 102.595 ;
        RECT 109.795 101.875 110.115 102.195 ;
        RECT 109.795 101.475 110.115 101.795 ;
        RECT 109.795 79.075 110.115 79.395 ;
        RECT 109.795 78.675 110.115 78.995 ;
        RECT 109.795 78.275 110.115 78.595 ;
        RECT 109.795 77.875 110.115 78.195 ;
        RECT 109.795 77.475 110.115 77.795 ;
        RECT 111.165 151.075 111.485 151.395 ;
        RECT 111.165 150.675 111.485 150.995 ;
        RECT 111.165 150.275 111.485 150.595 ;
        RECT 111.165 149.875 111.485 150.195 ;
        RECT 111.165 149.475 111.485 149.795 ;
        RECT 111.165 127.075 111.485 127.395 ;
        RECT 111.165 126.675 111.485 126.995 ;
        RECT 111.165 126.275 111.485 126.595 ;
        RECT 111.165 125.875 111.485 126.195 ;
        RECT 111.165 125.475 111.485 125.795 ;
        RECT 111.165 103.075 111.485 103.395 ;
        RECT 111.165 102.675 111.485 102.995 ;
        RECT 111.165 102.275 111.485 102.595 ;
        RECT 111.165 101.875 111.485 102.195 ;
        RECT 111.165 101.475 111.485 101.795 ;
        RECT 111.165 79.075 111.485 79.395 ;
        RECT 111.165 78.675 111.485 78.995 ;
        RECT 111.165 78.275 111.485 78.595 ;
        RECT 111.165 77.875 111.485 78.195 ;
        RECT 111.165 77.475 111.485 77.795 ;
        RECT 112.535 151.075 112.855 151.395 ;
        RECT 112.535 150.675 112.855 150.995 ;
        RECT 112.535 150.275 112.855 150.595 ;
        RECT 112.535 149.875 112.855 150.195 ;
        RECT 112.535 149.475 112.855 149.795 ;
        RECT 112.535 127.075 112.855 127.395 ;
        RECT 112.535 126.675 112.855 126.995 ;
        RECT 112.535 126.275 112.855 126.595 ;
        RECT 112.535 125.875 112.855 126.195 ;
        RECT 112.535 125.475 112.855 125.795 ;
        RECT 112.535 103.075 112.855 103.395 ;
        RECT 112.535 102.675 112.855 102.995 ;
        RECT 112.535 102.275 112.855 102.595 ;
        RECT 112.535 101.875 112.855 102.195 ;
        RECT 112.535 101.475 112.855 101.795 ;
        RECT 112.535 79.075 112.855 79.395 ;
        RECT 112.535 78.675 112.855 78.995 ;
        RECT 112.535 78.275 112.855 78.595 ;
        RECT 112.535 77.875 112.855 78.195 ;
        RECT 112.535 77.475 112.855 77.795 ;
        RECT 123.000 163.075 123.320 163.395 ;
        RECT 123.000 162.675 123.320 162.995 ;
        RECT 123.000 162.275 123.320 162.595 ;
        RECT 123.000 161.875 123.320 162.195 ;
        RECT 123.000 161.475 123.320 161.795 ;
        RECT 123.000 139.075 123.320 139.395 ;
        RECT 123.000 138.675 123.320 138.995 ;
        RECT 123.000 138.275 123.320 138.595 ;
        RECT 123.000 137.875 123.320 138.195 ;
        RECT 123.000 137.475 123.320 137.795 ;
        RECT 123.000 115.075 123.320 115.395 ;
        RECT 123.000 114.675 123.320 114.995 ;
        RECT 123.000 114.275 123.320 114.595 ;
        RECT 123.000 113.875 123.320 114.195 ;
        RECT 123.000 113.475 123.320 113.795 ;
        RECT 123.000 91.075 123.320 91.395 ;
        RECT 123.000 90.675 123.320 90.995 ;
        RECT 123.000 90.275 123.320 90.595 ;
        RECT 123.000 89.875 123.320 90.195 ;
        RECT 123.000 89.475 123.320 89.795 ;
        RECT 124.370 163.075 124.690 163.395 ;
        RECT 124.370 162.675 124.690 162.995 ;
        RECT 124.370 162.275 124.690 162.595 ;
        RECT 124.370 161.875 124.690 162.195 ;
        RECT 124.370 161.475 124.690 161.795 ;
        RECT 124.370 139.075 124.690 139.395 ;
        RECT 124.370 138.675 124.690 138.995 ;
        RECT 124.370 138.275 124.690 138.595 ;
        RECT 124.370 137.875 124.690 138.195 ;
        RECT 124.370 137.475 124.690 137.795 ;
        RECT 124.370 115.075 124.690 115.395 ;
        RECT 124.370 114.675 124.690 114.995 ;
        RECT 124.370 114.275 124.690 114.595 ;
        RECT 124.370 113.875 124.690 114.195 ;
        RECT 124.370 113.475 124.690 113.795 ;
        RECT 124.370 91.075 124.690 91.395 ;
        RECT 124.370 90.675 124.690 90.995 ;
        RECT 124.370 90.275 124.690 90.595 ;
        RECT 124.370 89.875 124.690 90.195 ;
        RECT 124.370 89.475 124.690 89.795 ;
        RECT 125.615 67.075 125.935 67.395 ;
        RECT 125.615 66.675 125.935 66.995 ;
        RECT 125.615 66.275 125.935 66.595 ;
        RECT 125.615 65.875 125.935 66.195 ;
        RECT 125.615 65.475 125.935 65.795 ;
        RECT 146.685 210.145 147.005 210.465 ;
        RECT 147.085 210.145 147.405 210.465 ;
        RECT 147.485 210.145 147.805 210.465 ;
        RECT 140.605 208.080 140.925 208.400 ;
        RECT 141.005 208.080 141.325 208.400 ;
        RECT 141.405 208.080 141.725 208.400 ;
        RECT 141.805 208.080 142.125 208.400 ;
        RECT 142.205 208.080 142.525 208.400 ;
        RECT 129.570 206.680 129.890 207.000 ;
        RECT 129.570 206.280 129.890 206.600 ;
        RECT 129.570 205.880 129.890 206.200 ;
        RECT 129.570 205.480 129.890 205.800 ;
        RECT 129.570 205.080 129.890 205.400 ;
        RECT 129.570 204.680 129.890 205.000 ;
        RECT 129.570 204.280 129.890 204.600 ;
        RECT 129.570 203.880 129.890 204.200 ;
        RECT 129.570 203.480 129.890 203.800 ;
        RECT 129.570 203.080 129.890 203.400 ;
        RECT 129.570 202.680 129.890 203.000 ;
        RECT 129.570 202.280 129.890 202.600 ;
        RECT 129.570 201.880 129.890 202.200 ;
        RECT 129.570 201.480 129.890 201.800 ;
        RECT 129.570 201.080 129.890 201.400 ;
        RECT 129.570 200.680 129.890 201.000 ;
        RECT 129.570 200.280 129.890 200.600 ;
        RECT 129.570 199.880 129.890 200.200 ;
        RECT 129.570 199.480 129.890 199.800 ;
        RECT 129.570 199.080 129.890 199.400 ;
        RECT 129.570 198.680 129.890 199.000 ;
        RECT 129.570 198.280 129.890 198.600 ;
        RECT 129.570 197.880 129.890 198.200 ;
        RECT 129.570 197.480 129.890 197.800 ;
        RECT 129.570 197.080 129.890 197.400 ;
        RECT 129.570 196.680 129.890 197.000 ;
        RECT 129.570 196.280 129.890 196.600 ;
        RECT 129.570 195.880 129.890 196.200 ;
        RECT 129.570 195.480 129.890 195.800 ;
        RECT 129.570 195.080 129.890 195.400 ;
        RECT 129.570 194.680 129.890 195.000 ;
        RECT 129.570 194.280 129.890 194.600 ;
        RECT 129.570 193.880 129.890 194.200 ;
        RECT 129.570 193.480 129.890 193.800 ;
        RECT 129.570 193.080 129.890 193.400 ;
        RECT 129.570 192.680 129.890 193.000 ;
        RECT 129.570 192.280 129.890 192.600 ;
        RECT 129.570 191.880 129.890 192.200 ;
        RECT 129.570 191.480 129.890 191.800 ;
        RECT 129.570 191.080 129.890 191.400 ;
        RECT 129.570 190.680 129.890 191.000 ;
        RECT 129.570 190.280 129.890 190.600 ;
        RECT 129.570 189.880 129.890 190.200 ;
        RECT 129.570 189.480 129.890 189.800 ;
        RECT 129.570 189.080 129.890 189.400 ;
        RECT 129.570 188.680 129.890 189.000 ;
        RECT 129.570 188.280 129.890 188.600 ;
        RECT 129.570 187.880 129.890 188.200 ;
        RECT 129.570 187.480 129.890 187.800 ;
        RECT 129.570 187.080 129.890 187.400 ;
        RECT 129.570 186.680 129.890 187.000 ;
        RECT 129.570 186.280 129.890 186.600 ;
        RECT 129.570 185.880 129.890 186.200 ;
        RECT 129.570 185.480 129.890 185.800 ;
        RECT 129.570 185.080 129.890 185.400 ;
        RECT 129.570 184.680 129.890 185.000 ;
        RECT 129.570 181.385 129.890 181.705 ;
        RECT 129.570 180.985 129.890 181.305 ;
        RECT 129.570 180.585 129.890 180.905 ;
        RECT 129.570 180.185 129.890 180.505 ;
        RECT 129.570 179.785 129.890 180.105 ;
        RECT 129.570 179.385 129.890 179.705 ;
        RECT 129.570 178.985 129.890 179.305 ;
        RECT 129.570 178.585 129.890 178.905 ;
        RECT 129.570 178.185 129.890 178.505 ;
        RECT 129.570 177.785 129.890 178.105 ;
        RECT 129.570 177.385 129.890 177.705 ;
        RECT 129.570 176.985 129.890 177.305 ;
        RECT 129.570 176.585 129.890 176.905 ;
        RECT 129.570 176.185 129.890 176.505 ;
        RECT 129.570 175.785 129.890 176.105 ;
        RECT 129.570 175.385 129.890 175.705 ;
        RECT 129.570 174.985 129.890 175.305 ;
        RECT 129.570 174.585 129.890 174.905 ;
        RECT 129.570 174.185 129.890 174.505 ;
        RECT 129.570 173.785 129.890 174.105 ;
        RECT 129.570 173.385 129.890 173.705 ;
        RECT 129.570 172.985 129.890 173.305 ;
        RECT 129.570 172.585 129.890 172.905 ;
        RECT 129.570 172.185 129.890 172.505 ;
        RECT 129.570 171.785 129.890 172.105 ;
        RECT 129.570 171.385 129.890 171.705 ;
        RECT 129.570 170.985 129.890 171.305 ;
        RECT 129.570 170.585 129.890 170.905 ;
        RECT 129.570 170.185 129.890 170.505 ;
        RECT 129.570 169.785 129.890 170.105 ;
        RECT 129.570 169.385 129.890 169.705 ;
        RECT 129.570 168.985 129.890 169.305 ;
        RECT 129.570 168.585 129.890 168.905 ;
        RECT 129.570 168.185 129.890 168.505 ;
        RECT 129.570 167.785 129.890 168.105 ;
        RECT 129.570 167.385 129.890 167.705 ;
        RECT 129.570 166.985 129.890 167.305 ;
        RECT 129.570 166.585 129.890 166.905 ;
        RECT 129.570 166.185 129.890 166.505 ;
        RECT 129.570 165.785 129.890 166.105 ;
        RECT 129.570 165.385 129.890 165.705 ;
        RECT 129.570 164.985 129.890 165.305 ;
        RECT 129.570 164.585 129.890 164.905 ;
        RECT 129.570 164.185 129.890 164.505 ;
        RECT 129.570 163.785 129.890 164.105 ;
        RECT 129.570 163.385 129.890 163.705 ;
        RECT 129.570 162.985 129.890 163.305 ;
        RECT 129.570 162.585 129.890 162.905 ;
        RECT 129.570 162.185 129.890 162.505 ;
        RECT 129.570 161.785 129.890 162.105 ;
        RECT 129.570 161.385 129.890 161.705 ;
        RECT 129.570 160.985 129.890 161.305 ;
        RECT 129.570 160.585 129.890 160.905 ;
        RECT 129.570 160.185 129.890 160.505 ;
        RECT 129.570 159.785 129.890 160.105 ;
        RECT 129.570 159.385 129.890 159.705 ;
        RECT 129.570 157.585 129.890 157.905 ;
        RECT 129.570 157.185 129.890 157.505 ;
        RECT 129.570 156.785 129.890 157.105 ;
        RECT 129.570 156.385 129.890 156.705 ;
        RECT 129.570 155.985 129.890 156.305 ;
        RECT 129.570 155.585 129.890 155.905 ;
        RECT 129.570 155.185 129.890 155.505 ;
        RECT 129.570 154.785 129.890 155.105 ;
        RECT 129.570 154.385 129.890 154.705 ;
        RECT 129.570 153.985 129.890 154.305 ;
        RECT 129.570 153.585 129.890 153.905 ;
        RECT 129.570 153.185 129.890 153.505 ;
        RECT 129.570 152.785 129.890 153.105 ;
        RECT 129.570 152.385 129.890 152.705 ;
        RECT 129.570 151.985 129.890 152.305 ;
        RECT 129.570 151.585 129.890 151.905 ;
        RECT 129.570 151.185 129.890 151.505 ;
        RECT 129.570 150.785 129.890 151.105 ;
        RECT 129.570 150.385 129.890 150.705 ;
        RECT 129.570 149.985 129.890 150.305 ;
        RECT 129.570 149.585 129.890 149.905 ;
        RECT 129.570 149.185 129.890 149.505 ;
        RECT 129.570 148.785 129.890 149.105 ;
        RECT 129.570 148.385 129.890 148.705 ;
        RECT 129.570 147.985 129.890 148.305 ;
        RECT 129.570 147.585 129.890 147.905 ;
        RECT 129.570 147.185 129.890 147.505 ;
        RECT 129.570 146.785 129.890 147.105 ;
        RECT 129.570 146.385 129.890 146.705 ;
        RECT 129.570 145.985 129.890 146.305 ;
        RECT 129.570 145.585 129.890 145.905 ;
        RECT 129.570 145.185 129.890 145.505 ;
        RECT 129.570 144.785 129.890 145.105 ;
        RECT 129.570 144.385 129.890 144.705 ;
        RECT 129.570 143.985 129.890 144.305 ;
        RECT 129.570 143.585 129.890 143.905 ;
        RECT 129.570 143.185 129.890 143.505 ;
        RECT 129.570 142.785 129.890 143.105 ;
        RECT 129.570 142.385 129.890 142.705 ;
        RECT 129.570 141.985 129.890 142.305 ;
        RECT 129.570 141.585 129.890 141.905 ;
        RECT 129.570 141.185 129.890 141.505 ;
        RECT 129.570 140.785 129.890 141.105 ;
        RECT 129.570 140.385 129.890 140.705 ;
        RECT 129.570 139.985 129.890 140.305 ;
        RECT 129.570 139.585 129.890 139.905 ;
        RECT 129.570 139.185 129.890 139.505 ;
        RECT 129.570 138.785 129.890 139.105 ;
        RECT 129.570 138.385 129.890 138.705 ;
        RECT 129.570 137.985 129.890 138.305 ;
        RECT 129.570 137.585 129.890 137.905 ;
        RECT 129.570 137.185 129.890 137.505 ;
        RECT 129.570 136.785 129.890 137.105 ;
        RECT 129.570 136.385 129.890 136.705 ;
        RECT 129.570 135.985 129.890 136.305 ;
        RECT 129.570 135.585 129.890 135.905 ;
        RECT 129.570 133.785 129.890 134.105 ;
        RECT 129.570 133.385 129.890 133.705 ;
        RECT 129.570 132.985 129.890 133.305 ;
        RECT 129.570 132.585 129.890 132.905 ;
        RECT 129.570 132.185 129.890 132.505 ;
        RECT 129.570 131.785 129.890 132.105 ;
        RECT 129.570 131.385 129.890 131.705 ;
        RECT 129.570 130.985 129.890 131.305 ;
        RECT 129.570 130.585 129.890 130.905 ;
        RECT 129.570 130.185 129.890 130.505 ;
        RECT 129.570 129.785 129.890 130.105 ;
        RECT 129.570 129.385 129.890 129.705 ;
        RECT 129.570 128.985 129.890 129.305 ;
        RECT 129.570 128.585 129.890 128.905 ;
        RECT 129.570 128.185 129.890 128.505 ;
        RECT 129.570 127.785 129.890 128.105 ;
        RECT 129.570 127.385 129.890 127.705 ;
        RECT 129.570 126.985 129.890 127.305 ;
        RECT 129.570 126.585 129.890 126.905 ;
        RECT 129.570 126.185 129.890 126.505 ;
        RECT 129.570 125.785 129.890 126.105 ;
        RECT 129.570 125.385 129.890 125.705 ;
        RECT 129.570 124.985 129.890 125.305 ;
        RECT 129.570 124.585 129.890 124.905 ;
        RECT 129.570 124.185 129.890 124.505 ;
        RECT 129.570 123.785 129.890 124.105 ;
        RECT 129.570 123.385 129.890 123.705 ;
        RECT 129.570 122.985 129.890 123.305 ;
        RECT 129.570 122.585 129.890 122.905 ;
        RECT 129.570 122.185 129.890 122.505 ;
        RECT 129.570 121.785 129.890 122.105 ;
        RECT 129.570 121.385 129.890 121.705 ;
        RECT 129.570 120.985 129.890 121.305 ;
        RECT 129.570 120.585 129.890 120.905 ;
        RECT 129.570 120.185 129.890 120.505 ;
        RECT 129.570 119.785 129.890 120.105 ;
        RECT 129.570 119.385 129.890 119.705 ;
        RECT 129.570 118.985 129.890 119.305 ;
        RECT 129.570 118.585 129.890 118.905 ;
        RECT 129.570 118.185 129.890 118.505 ;
        RECT 129.570 117.785 129.890 118.105 ;
        RECT 129.570 117.385 129.890 117.705 ;
        RECT 129.570 116.985 129.890 117.305 ;
        RECT 129.570 116.585 129.890 116.905 ;
        RECT 129.570 116.185 129.890 116.505 ;
        RECT 129.570 115.785 129.890 116.105 ;
        RECT 129.570 115.385 129.890 115.705 ;
        RECT 129.570 114.985 129.890 115.305 ;
        RECT 129.570 114.585 129.890 114.905 ;
        RECT 129.570 114.185 129.890 114.505 ;
        RECT 129.570 113.785 129.890 114.105 ;
        RECT 129.570 113.385 129.890 113.705 ;
        RECT 129.570 112.985 129.890 113.305 ;
        RECT 129.570 112.585 129.890 112.905 ;
        RECT 129.570 112.185 129.890 112.505 ;
        RECT 129.570 111.785 129.890 112.105 ;
        RECT 129.570 109.985 129.890 110.305 ;
        RECT 129.570 109.585 129.890 109.905 ;
        RECT 129.570 109.185 129.890 109.505 ;
        RECT 129.570 108.785 129.890 109.105 ;
        RECT 129.570 108.385 129.890 108.705 ;
        RECT 129.570 107.985 129.890 108.305 ;
        RECT 129.570 107.585 129.890 107.905 ;
        RECT 129.570 107.185 129.890 107.505 ;
        RECT 129.570 106.785 129.890 107.105 ;
        RECT 129.570 106.385 129.890 106.705 ;
        RECT 129.570 105.985 129.890 106.305 ;
        RECT 129.570 105.585 129.890 105.905 ;
        RECT 129.570 105.185 129.890 105.505 ;
        RECT 129.570 104.785 129.890 105.105 ;
        RECT 129.570 104.385 129.890 104.705 ;
        RECT 129.570 103.985 129.890 104.305 ;
        RECT 129.570 103.585 129.890 103.905 ;
        RECT 129.570 103.185 129.890 103.505 ;
        RECT 129.570 102.785 129.890 103.105 ;
        RECT 129.570 102.385 129.890 102.705 ;
        RECT 129.570 101.985 129.890 102.305 ;
        RECT 129.570 101.585 129.890 101.905 ;
        RECT 129.570 101.185 129.890 101.505 ;
        RECT 129.570 100.785 129.890 101.105 ;
        RECT 129.570 100.385 129.890 100.705 ;
        RECT 129.570 99.985 129.890 100.305 ;
        RECT 129.570 99.585 129.890 99.905 ;
        RECT 129.570 99.185 129.890 99.505 ;
        RECT 129.570 98.785 129.890 99.105 ;
        RECT 129.570 98.385 129.890 98.705 ;
        RECT 129.570 97.985 129.890 98.305 ;
        RECT 129.570 97.585 129.890 97.905 ;
        RECT 129.570 97.185 129.890 97.505 ;
        RECT 129.570 96.785 129.890 97.105 ;
        RECT 129.570 96.385 129.890 96.705 ;
        RECT 129.570 95.985 129.890 96.305 ;
        RECT 129.570 95.585 129.890 95.905 ;
        RECT 129.570 95.185 129.890 95.505 ;
        RECT 129.570 94.785 129.890 95.105 ;
        RECT 129.570 94.385 129.890 94.705 ;
        RECT 129.570 93.985 129.890 94.305 ;
        RECT 129.570 93.585 129.890 93.905 ;
        RECT 129.570 93.185 129.890 93.505 ;
        RECT 129.570 92.785 129.890 93.105 ;
        RECT 129.570 92.385 129.890 92.705 ;
        RECT 129.570 91.985 129.890 92.305 ;
        RECT 129.570 91.585 129.890 91.905 ;
        RECT 129.570 91.185 129.890 91.505 ;
        RECT 129.570 90.785 129.890 91.105 ;
        RECT 129.570 90.385 129.890 90.705 ;
        RECT 129.570 89.985 129.890 90.305 ;
        RECT 129.570 89.585 129.890 89.905 ;
        RECT 129.570 89.185 129.890 89.505 ;
        RECT 129.570 88.785 129.890 89.105 ;
        RECT 129.570 88.385 129.890 88.705 ;
        RECT 129.570 87.985 129.890 88.305 ;
        RECT 129.570 86.185 129.890 86.505 ;
        RECT 129.570 85.785 129.890 86.105 ;
        RECT 129.570 85.385 129.890 85.705 ;
        RECT 129.570 84.985 129.890 85.305 ;
        RECT 129.570 84.585 129.890 84.905 ;
        RECT 129.570 84.185 129.890 84.505 ;
        RECT 129.570 83.785 129.890 84.105 ;
        RECT 129.570 83.385 129.890 83.705 ;
        RECT 129.570 82.985 129.890 83.305 ;
        RECT 129.570 82.585 129.890 82.905 ;
        RECT 129.570 82.185 129.890 82.505 ;
        RECT 129.570 81.785 129.890 82.105 ;
        RECT 129.570 81.385 129.890 81.705 ;
        RECT 129.570 80.985 129.890 81.305 ;
        RECT 129.570 80.585 129.890 80.905 ;
        RECT 129.570 80.185 129.890 80.505 ;
        RECT 129.570 79.785 129.890 80.105 ;
        RECT 129.570 79.385 129.890 79.705 ;
        RECT 129.570 78.985 129.890 79.305 ;
        RECT 129.570 78.585 129.890 78.905 ;
        RECT 129.570 78.185 129.890 78.505 ;
        RECT 129.570 77.785 129.890 78.105 ;
        RECT 129.570 77.385 129.890 77.705 ;
        RECT 129.570 76.985 129.890 77.305 ;
        RECT 129.570 76.585 129.890 76.905 ;
        RECT 129.570 76.185 129.890 76.505 ;
        RECT 129.570 75.785 129.890 76.105 ;
        RECT 129.570 75.385 129.890 75.705 ;
        RECT 129.570 74.985 129.890 75.305 ;
        RECT 129.570 74.585 129.890 74.905 ;
        RECT 129.570 74.185 129.890 74.505 ;
        RECT 129.570 73.785 129.890 74.105 ;
        RECT 129.570 73.385 129.890 73.705 ;
        RECT 129.570 72.985 129.890 73.305 ;
        RECT 129.570 72.585 129.890 72.905 ;
        RECT 129.570 72.185 129.890 72.505 ;
        RECT 129.570 71.785 129.890 72.105 ;
        RECT 129.570 71.385 129.890 71.705 ;
        RECT 129.570 70.985 129.890 71.305 ;
        RECT 129.570 70.585 129.890 70.905 ;
        RECT 129.570 70.185 129.890 70.505 ;
        RECT 129.570 69.785 129.890 70.105 ;
        RECT 129.570 69.385 129.890 69.705 ;
        RECT 129.570 68.985 129.890 69.305 ;
        RECT 129.570 68.585 129.890 68.905 ;
        RECT 129.570 68.185 129.890 68.505 ;
        RECT 129.570 67.785 129.890 68.105 ;
        RECT 129.570 67.385 129.890 67.705 ;
        RECT 129.570 66.985 129.890 67.305 ;
        RECT 129.570 66.585 129.890 66.905 ;
        RECT 129.570 66.185 129.890 66.505 ;
        RECT 129.570 65.785 129.890 66.105 ;
        RECT 129.570 65.385 129.890 65.705 ;
        RECT 129.570 64.985 129.890 65.305 ;
        RECT 129.570 64.585 129.890 64.905 ;
        RECT 129.570 64.185 129.890 64.505 ;
        RECT 129.570 62.385 129.890 62.705 ;
        RECT 129.570 61.985 129.890 62.305 ;
        RECT 129.570 61.585 129.890 61.905 ;
        RECT 129.570 61.185 129.890 61.505 ;
        RECT 129.570 60.785 129.890 61.105 ;
        RECT 129.570 60.385 129.890 60.705 ;
        RECT 129.570 59.985 129.890 60.305 ;
        RECT 129.570 59.585 129.890 59.905 ;
        RECT 129.570 59.185 129.890 59.505 ;
        RECT 129.570 58.785 129.890 59.105 ;
        RECT 129.570 58.385 129.890 58.705 ;
        RECT 129.570 57.985 129.890 58.305 ;
        RECT 129.570 57.585 129.890 57.905 ;
        RECT 129.570 57.185 129.890 57.505 ;
        RECT 129.570 56.785 129.890 57.105 ;
        RECT 129.570 56.385 129.890 56.705 ;
        RECT 129.570 55.985 129.890 56.305 ;
        RECT 129.570 55.585 129.890 55.905 ;
        RECT 129.570 55.185 129.890 55.505 ;
        RECT 129.570 54.785 129.890 55.105 ;
        RECT 129.570 54.385 129.890 54.705 ;
        RECT 129.570 53.985 129.890 54.305 ;
        RECT 129.570 53.585 129.890 53.905 ;
        RECT 129.570 53.185 129.890 53.505 ;
        RECT 129.570 52.785 129.890 53.105 ;
        RECT 129.570 52.385 129.890 52.705 ;
        RECT 129.570 51.985 129.890 52.305 ;
        RECT 129.570 51.585 129.890 51.905 ;
        RECT 129.570 51.185 129.890 51.505 ;
        RECT 129.570 50.785 129.890 51.105 ;
        RECT 129.570 50.385 129.890 50.705 ;
        RECT 129.570 49.985 129.890 50.305 ;
        RECT 129.570 49.585 129.890 49.905 ;
        RECT 129.570 49.185 129.890 49.505 ;
        RECT 129.570 48.785 129.890 49.105 ;
        RECT 129.570 48.385 129.890 48.705 ;
        RECT 129.570 47.985 129.890 48.305 ;
        RECT 129.570 47.585 129.890 47.905 ;
        RECT 129.570 47.185 129.890 47.505 ;
        RECT 129.570 46.785 129.890 47.105 ;
        RECT 129.570 46.385 129.890 46.705 ;
        RECT 129.570 45.985 129.890 46.305 ;
        RECT 129.570 45.585 129.890 45.905 ;
        RECT 129.570 45.185 129.890 45.505 ;
        RECT 129.570 44.785 129.890 45.105 ;
        RECT 129.570 44.385 129.890 44.705 ;
        RECT 129.570 43.985 129.890 44.305 ;
        RECT 129.570 43.585 129.890 43.905 ;
        RECT 129.570 43.185 129.890 43.505 ;
        RECT 129.570 42.785 129.890 43.105 ;
        RECT 129.570 42.385 129.890 42.705 ;
        RECT 129.570 41.985 129.890 42.305 ;
        RECT 129.570 41.585 129.890 41.905 ;
        RECT 129.570 41.185 129.890 41.505 ;
        RECT 129.570 40.785 129.890 41.105 ;
        RECT 129.570 40.385 129.890 40.705 ;
        RECT 140.605 38.845 140.925 39.165 ;
        RECT 141.005 38.845 141.325 39.165 ;
        RECT 141.405 38.845 141.725 39.165 ;
        RECT 141.805 38.845 142.125 39.165 ;
        RECT 142.205 38.845 142.525 39.165 ;
        RECT 129.570 37.085 129.890 37.405 ;
        RECT 129.570 36.685 129.890 37.005 ;
        RECT 129.570 36.285 129.890 36.605 ;
        RECT 129.570 35.885 129.890 36.205 ;
        RECT 129.570 35.485 129.890 35.805 ;
        RECT 129.570 35.085 129.890 35.405 ;
        RECT 129.570 34.685 129.890 35.005 ;
        RECT 129.570 34.285 129.890 34.605 ;
        RECT 129.570 33.885 129.890 34.205 ;
        RECT 129.570 33.485 129.890 33.805 ;
        RECT 129.570 33.085 129.890 33.405 ;
        RECT 129.570 32.685 129.890 33.005 ;
        RECT 129.570 32.285 129.890 32.605 ;
        RECT 129.570 31.885 129.890 32.205 ;
        RECT 129.570 31.485 129.890 31.805 ;
        RECT 129.570 31.085 129.890 31.405 ;
        RECT 129.570 30.685 129.890 31.005 ;
        RECT 129.570 30.285 129.890 30.605 ;
        RECT 129.570 29.885 129.890 30.205 ;
        RECT 129.570 29.485 129.890 29.805 ;
        RECT 129.570 29.085 129.890 29.405 ;
        RECT 129.570 28.685 129.890 29.005 ;
        RECT 129.570 28.285 129.890 28.605 ;
        RECT 129.570 27.885 129.890 28.205 ;
        RECT 129.570 27.485 129.890 27.805 ;
        RECT 129.570 27.085 129.890 27.405 ;
        RECT 129.570 26.685 129.890 27.005 ;
        RECT 129.570 26.285 129.890 26.605 ;
        RECT 129.570 25.885 129.890 26.205 ;
        RECT 129.570 25.485 129.890 25.805 ;
        RECT 129.570 25.085 129.890 25.405 ;
        RECT 129.570 24.685 129.890 25.005 ;
        RECT 129.570 24.285 129.890 24.605 ;
        RECT 129.570 23.885 129.890 24.205 ;
        RECT 129.570 23.485 129.890 23.805 ;
        RECT 129.570 23.085 129.890 23.405 ;
        RECT 129.570 22.685 129.890 23.005 ;
        RECT 129.570 22.285 129.890 22.605 ;
        RECT 129.570 21.885 129.890 22.205 ;
        RECT 129.570 21.485 129.890 21.805 ;
        RECT 129.570 21.085 129.890 21.405 ;
        RECT 129.570 20.685 129.890 21.005 ;
        RECT 129.570 20.285 129.890 20.605 ;
        RECT 129.570 19.885 129.890 20.205 ;
        RECT 129.570 19.485 129.890 19.805 ;
        RECT 129.570 19.085 129.890 19.405 ;
        RECT 129.570 18.685 129.890 19.005 ;
        RECT 129.570 18.285 129.890 18.605 ;
        RECT 129.570 17.885 129.890 18.205 ;
        RECT 129.570 17.485 129.890 17.805 ;
        RECT 129.570 17.085 129.890 17.405 ;
        RECT 129.570 16.685 129.890 17.005 ;
        RECT 129.570 16.285 129.890 16.605 ;
        RECT 129.570 15.885 129.890 16.205 ;
        RECT 129.570 15.485 129.890 15.805 ;
        RECT 129.570 15.085 129.890 15.405 ;
        RECT 140.605 13.685 140.925 14.005 ;
        RECT 141.005 13.685 141.325 14.005 ;
        RECT 141.405 13.685 141.725 14.005 ;
        RECT 141.805 13.685 142.125 14.005 ;
        RECT 142.205 13.685 142.525 14.005 ;
        RECT 111.875 7.635 112.195 7.955 ;
        RECT 112.275 7.635 112.595 7.955 ;
        RECT 112.675 7.635 112.995 7.955 ;
        RECT 89.795 6.535 90.115 6.855 ;
        RECT 90.195 6.535 90.515 6.855 ;
        RECT 90.595 6.535 90.915 6.855 ;
        RECT 134.485 4.215 134.805 4.535 ;
        RECT 134.885 4.215 135.205 4.535 ;
        RECT 135.285 4.215 135.605 4.535 ;
        RECT 135.685 4.215 136.005 4.535 ;
        RECT 90.460 3.420 90.780 3.740 ;
        RECT 90.460 3.020 90.780 3.340 ;
        RECT 90.460 2.620 90.780 2.940 ;
        RECT 90.460 2.220 90.780 2.540 ;
        RECT 90.460 1.820 90.780 2.140 ;
        RECT 112.540 3.420 112.860 3.740 ;
        RECT 112.540 3.020 112.860 3.340 ;
        RECT 112.540 2.620 112.860 2.940 ;
        RECT 112.540 2.220 112.860 2.540 ;
        RECT 112.540 1.820 112.860 2.140 ;
        RECT 134.620 3.420 134.940 3.740 ;
        RECT 134.620 3.020 134.940 3.340 ;
        RECT 134.620 2.620 134.940 2.940 ;
        RECT 134.620 2.220 134.940 2.540 ;
        RECT 134.620 1.820 134.940 2.140 ;
        RECT 156.705 3.420 157.025 3.740 ;
        RECT 156.705 3.020 157.025 3.340 ;
        RECT 156.705 2.620 157.025 2.940 ;
        RECT 156.705 2.220 157.025 2.540 ;
        RECT 156.705 1.820 157.025 2.140 ;
      LAYER met4 ;
        RECT 3.990 220.760 4.290 225.760 ;
        RECT 7.670 220.760 7.970 225.760 ;
        RECT 11.350 220.760 11.650 225.760 ;
        RECT 15.030 220.760 15.330 225.760 ;
        RECT 18.710 220.760 19.010 225.760 ;
        RECT 22.390 220.760 22.690 225.760 ;
        RECT 26.070 220.760 26.370 225.760 ;
        RECT 29.750 220.760 30.050 225.760 ;
        RECT 33.430 220.760 33.730 225.760 ;
        RECT 37.110 220.760 37.410 225.760 ;
        RECT 40.790 220.760 41.090 225.760 ;
        RECT 44.470 220.760 44.770 225.760 ;
        RECT 48.150 220.760 48.450 225.760 ;
        RECT 51.830 220.760 52.130 225.760 ;
        RECT 55.510 220.760 55.810 225.760 ;
        RECT 59.190 220.760 59.490 225.760 ;
        RECT 62.870 220.760 63.170 225.760 ;
        RECT 66.550 220.760 66.850 225.760 ;
        RECT 70.230 220.760 70.530 225.760 ;
        RECT 73.910 220.760 74.210 225.760 ;
        RECT 77.590 220.760 77.890 225.760 ;
        RECT 81.270 220.760 81.570 225.760 ;
        RECT 1.000 5.000 2.500 220.760 ;
        RECT 3.975 219.260 4.305 220.760 ;
        RECT 7.655 219.260 7.985 220.760 ;
        RECT 11.335 219.260 11.665 220.760 ;
        RECT 15.015 219.260 15.345 220.760 ;
        RECT 18.695 219.260 19.025 220.760 ;
        RECT 22.375 219.260 22.705 220.760 ;
        RECT 26.055 219.260 26.385 220.760 ;
        RECT 29.735 219.260 30.065 220.760 ;
        RECT 33.415 219.260 33.745 220.760 ;
        RECT 37.095 219.260 37.425 220.760 ;
        RECT 40.775 219.260 41.105 220.760 ;
        RECT 44.455 219.260 44.785 220.760 ;
        RECT 48.135 219.260 48.465 220.760 ;
        RECT 49.000 163.435 50.500 220.760 ;
        RECT 51.815 219.260 52.145 220.760 ;
        RECT 55.495 219.260 55.825 220.760 ;
        RECT 59.175 219.260 59.505 220.760 ;
        RECT 62.855 219.260 63.185 220.760 ;
        RECT 66.535 219.260 66.865 220.760 ;
        RECT 70.215 219.260 70.545 220.760 ;
        RECT 73.895 219.260 74.225 220.760 ;
        RECT 77.575 219.260 77.905 220.760 ;
        RECT 81.255 219.260 81.585 220.760 ;
        RECT 84.950 174.845 85.250 225.760 ;
        RECT 84.935 173.715 85.265 174.845 ;
        RECT 88.630 173.745 88.930 225.760 ;
        RECT 92.310 224.760 92.610 225.760 ;
        RECT 95.990 224.760 96.290 225.760 ;
        RECT 99.670 224.760 99.970 225.760 ;
        RECT 103.350 224.760 103.650 225.760 ;
        RECT 107.030 224.760 107.330 225.760 ;
        RECT 110.710 224.760 111.010 225.760 ;
        RECT 114.390 224.760 114.690 225.760 ;
        RECT 118.070 224.760 118.370 225.760 ;
        RECT 121.750 224.760 122.050 225.760 ;
        RECT 125.430 224.760 125.730 225.760 ;
        RECT 129.110 224.760 129.410 225.760 ;
        RECT 132.790 224.760 133.090 225.760 ;
        RECT 136.470 224.760 136.770 225.760 ;
        RECT 140.150 224.760 140.450 225.760 ;
        RECT 143.830 225.650 144.130 225.760 ;
        RECT 143.830 224.760 144.135 225.650 ;
        RECT 143.835 212.130 144.135 224.760 ;
        RECT 143.005 211.800 144.135 212.130 ;
        RECT 147.510 210.470 147.810 225.760 ;
        RECT 151.190 224.760 151.490 225.760 ;
        RECT 154.870 224.760 155.170 225.760 ;
        RECT 158.550 224.760 158.850 225.760 ;
        RECT 146.680 210.140 147.810 210.470 ;
        RECT 140.600 207.940 142.530 208.540 ;
        RECT 88.615 172.615 88.945 173.745 ;
        RECT 129.470 163.435 130.070 207.140 ;
        RECT 141.930 206.745 142.530 207.940 ;
        RECT 131.325 184.935 153.135 206.745 ;
        RECT 141.930 184.775 142.530 184.935 ;
        RECT 141.930 181.450 142.530 181.520 ;
        RECT 49.000 161.435 130.070 163.435 ;
        RECT 49.000 139.435 50.500 161.435 ;
        RECT 52.500 149.435 127.725 151.435 ;
        RECT 129.470 139.435 130.070 161.435 ;
        RECT 131.325 159.640 153.135 181.450 ;
        RECT 141.930 157.650 142.530 159.640 ;
        RECT 49.000 137.435 130.070 139.435 ;
        RECT 49.000 115.435 50.500 137.435 ;
        RECT 52.500 125.435 127.725 127.435 ;
        RECT 129.470 115.435 130.070 137.435 ;
        RECT 131.325 135.840 153.135 157.650 ;
        RECT 141.930 133.850 142.530 135.840 ;
        RECT 49.000 113.435 130.070 115.435 ;
        RECT 49.000 91.435 50.500 113.435 ;
        RECT 52.500 101.435 127.725 103.435 ;
        RECT 129.470 91.435 130.070 113.435 ;
        RECT 131.325 112.040 153.135 133.850 ;
        RECT 141.930 110.050 142.530 112.040 ;
        RECT 49.000 89.435 130.070 91.435 ;
        RECT 49.000 67.435 50.500 89.435 ;
        RECT 71.350 81.860 87.210 82.860 ;
        RECT 52.500 77.435 127.725 79.435 ;
        RECT 129.470 67.435 130.070 89.435 ;
        RECT 131.325 88.240 153.135 110.050 ;
        RECT 141.930 86.250 142.530 88.240 ;
        RECT 49.000 65.435 130.070 67.435 ;
        RECT 49.000 5.000 50.500 65.435 ;
        RECT 129.470 14.945 130.070 65.435 ;
        RECT 131.325 64.440 153.135 86.250 ;
        RECT 141.930 62.450 142.530 64.440 ;
        RECT 131.325 40.640 153.135 62.450 ;
        RECT 141.930 39.305 142.530 40.640 ;
        RECT 140.600 38.705 142.530 39.305 ;
        RECT 141.930 37.150 142.530 37.345 ;
        RECT 131.325 15.340 153.135 37.150 ;
        RECT 141.930 14.145 142.530 15.340 ;
        RECT 140.600 13.545 142.530 14.145 ;
        RECT 111.870 7.495 113.000 8.095 ;
        RECT 89.790 6.395 90.920 6.995 ;
        RECT 2.000 0.000 2.600 1.000 ;
        RECT 24.080 0.000 24.680 1.000 ;
        RECT 46.160 0.000 46.760 1.000 ;
        RECT 68.240 0.000 68.840 1.000 ;
        RECT 90.320 0.000 90.920 6.395 ;
        RECT 112.400 0.000 113.000 7.495 ;
        RECT 134.480 4.075 136.010 4.675 ;
        RECT 134.480 0.000 135.080 4.075 ;
        RECT 156.565 1.000 157.165 3.750 ;
        RECT 156.560 0.345 157.165 1.000 ;
        RECT 156.560 0.000 157.160 0.345 ;
  END
END tt_um_lcasimon_Tdc
END LIBRARY

