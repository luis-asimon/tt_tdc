MACRO System
  CLASS BLOCK ;
  FOREIGN System ;
  ORIGIN 18.005 48.000 ;
  SIZE 225.305 BY 157.265 ;
  PIN CL
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER met3 ;
        RECT 189.045 18.205 189.645 18.805 ;
    END
  END CL
  PIN Vout
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER met3 ;
        RECT 189.045 27.225 189.645 27.825 ;
    END
  END Vout
  PIN VoutN
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER met3 ;
        RECT 189.045 34.665 189.645 35.265 ;
    END
  END VoutN
  PIN CH
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER met3 ;
        RECT 189.045 41.985 189.645 42.585 ;
    END
  END CH
  PIN Vcap
    ANTENNAGATEAREA 32.000000 ;
    ANTENNADIFFAREA 1.960000 ;
    PORT
      LAYER met3 ;
        RECT 189.005 75.640 189.605 76.240 ;
    END
  END Vcap
  PIN VL
    ANTENNAGATEAREA 16.000000 ;
    ANTENNADIFFAREA 1.344000 ;
    PORT
      LAYER met3 ;
        RECT 189.315 68.715 189.645 69.045 ;
    END
  END VL
  PIN VH
    ANTENNAGATEAREA 16.000000 ;
    ANTENNADIFFAREA 1.344000 ;
    PORT
      LAYER met3 ;
        RECT 0.605 68.715 0.935 69.045 ;
    END
  END VH
  PIN VSS
    ANTENNAGATEAREA 77.360001 ;
    ANTENNADIFFAREA 179.072891 ;
    PORT
      LAYER met3 ;
        RECT 44.215 0.000 47.215 3.000 ;
    END
  END VSS
  PIN VDD
    ANTENNAGATEAREA 124.879997 ;
    ANTENNADIFFAREA 204.406494 ;
    PORT
      LAYER met3 ;
        RECT 44.215 3.500 47.215 6.500 ;
    END
  END VDD
  PIN ResetCH
    ANTENNAGATEAREA 1.200000 ;
    PORT
      LAYER met3 ;
        RECT 0.605 71.355 0.935 71.685 ;
    END
  END ResetCH
  PIN Reset
    ANTENNAGATEAREA 0.420000 ;
    PORT
      LAYER met3 ;
        RECT 189.275 78.395 189.605 78.725 ;
    END
  END Reset
  PIN Pulse
    ANTENNAGATEAREA 2.220000 ;
    PORT
      LAYER met3 ;
        RECT 0.605 66.375 0.935 66.705 ;
    END
  END Pulse
  PIN Iin
    ANTENNAGATEAREA 86.799995 ;
    ANTENNADIFFAREA 3.136000 ;
    PORT
      LAYER met3 ;
        RECT 0.600 74.680 0.930 75.010 ;
    END
  END Iin
  OBS
      LAYER pwell ;
        RECT 137.040 77.795 147.330 78.225 ;
        RECT 42.640 76.550 130.970 76.980 ;
        RECT 42.640 73.140 43.070 76.550 ;
        RECT 43.230 75.050 130.380 76.010 ;
        RECT 43.230 73.680 130.380 74.640 ;
        RECT 130.540 73.140 130.970 76.550 ;
        RECT 137.040 75.755 137.470 77.795 ;
        RECT 137.630 76.295 146.740 77.255 ;
        RECT 146.900 75.755 147.330 77.795 ;
        RECT 137.040 75.325 147.330 75.755 ;
        RECT 42.640 72.710 130.970 73.140 ;
        RECT 89.430 71.835 98.000 72.710 ;
        RECT 89.430 69.495 89.860 71.835 ;
        RECT 90.020 70.035 97.410 71.295 ;
        RECT 97.570 69.495 98.000 71.835 ;
        RECT 89.430 69.065 98.000 69.495 ;
        RECT 123.630 72.265 130.970 72.710 ;
        RECT 123.630 71.835 132.200 72.265 ;
        RECT 123.630 69.495 124.060 71.835 ;
        RECT 124.220 70.035 131.610 71.295 ;
        RECT 131.770 69.495 132.200 71.835 ;
        RECT 123.630 69.065 132.200 69.495 ;
        RECT 89.430 68.695 93.465 69.065 ;
        RECT 89.195 68.265 93.465 68.695 ;
        RECT 89.195 66.225 89.625 68.265 ;
        RECT 89.785 66.765 92.875 67.725 ;
        RECT 93.035 66.225 93.465 68.265 ;
        RECT 89.195 65.795 93.465 66.225 ;
      LAYER nwell ;
        RECT 33.400 61.395 38.710 65.355 ;
        RECT 93.775 65.195 98.225 68.745 ;
      LAYER pwell ;
        RECT 123.630 68.695 127.665 69.065 ;
      LAYER nwell ;
        RECT 136.950 68.745 142.260 75.005 ;
      LAYER pwell ;
        RECT 142.290 74.955 147.330 75.325 ;
        RECT 142.290 74.525 147.420 74.955 ;
        RECT 142.290 69.770 142.720 74.525 ;
        RECT 142.880 73.025 146.830 73.985 ;
        RECT 142.880 70.310 146.830 71.270 ;
        RECT 146.990 69.770 147.420 74.525 ;
        RECT 142.290 69.340 147.420 69.770 ;
        RECT 123.395 68.265 127.665 68.695 ;
        RECT 123.395 66.225 123.825 68.265 ;
        RECT 123.985 66.765 127.075 67.725 ;
        RECT 127.235 66.225 127.665 68.265 ;
        RECT 123.395 65.795 127.665 66.225 ;
      LAYER nwell ;
        RECT 127.975 65.590 147.660 68.745 ;
        RECT 127.975 65.195 144.740 65.590 ;
      LAYER pwell ;
        RECT 33.450 58.890 33.880 61.295 ;
        RECT 34.080 59.065 38.030 60.325 ;
        RECT 38.230 58.890 38.660 61.295 ;
      LAYER nwell ;
        RECT 42.550 59.455 144.740 65.195 ;
      LAYER pwell ;
        RECT 33.450 58.460 38.660 58.890 ;
      LAYER nwell ;
        RECT 55.800 46.900 95.830 53.790 ;
        RECT 93.960 46.285 95.830 46.900 ;
      LAYER pwell ;
        RECT 55.850 45.055 65.300 45.485 ;
        RECT 55.850 43.215 56.280 45.055 ;
        RECT 56.480 43.755 64.670 44.515 ;
        RECT 64.870 43.215 65.300 45.055 ;
        RECT 55.850 42.785 65.300 43.215 ;
        RECT 69.060 45.055 90.190 45.485 ;
        RECT 69.060 43.215 69.490 45.055 ;
        RECT 69.690 43.755 89.560 44.515 ;
        RECT 89.760 43.215 90.190 45.055 ;
        RECT 69.060 42.785 90.190 43.215 ;
      LAYER nwell ;
        RECT 93.960 42.325 118.630 46.285 ;
        RECT 124.280 42.310 129.590 46.270 ;
        RECT 134.940 42.310 144.550 46.270 ;
        RECT 69.010 38.480 90.240 41.780 ;
      LAYER pwell ;
        RECT 94.010 39.845 94.440 42.250 ;
        RECT 94.640 40.045 117.950 40.805 ;
        RECT 118.150 39.845 118.580 42.250 ;
        RECT 94.010 39.415 118.580 39.845 ;
        RECT 124.330 39.805 124.760 42.210 ;
        RECT 124.960 39.980 128.910 41.240 ;
        RECT 129.110 39.805 129.540 42.210 ;
        RECT 124.330 39.375 129.540 39.805 ;
        RECT 134.990 39.805 135.420 42.210 ;
        RECT 135.620 39.980 143.870 41.240 ;
        RECT 144.070 39.805 144.500 42.210 ;
        RECT 134.990 39.375 144.500 39.805 ;
        RECT 124.680 37.785 129.890 38.215 ;
        RECT 64.570 36.900 94.740 37.330 ;
        RECT 64.570 32.320 65.000 36.900 ;
        RECT 65.160 35.600 94.150 36.360 ;
        RECT 65.560 32.860 93.750 33.620 ;
        RECT 94.310 32.320 94.740 36.900 ;
        RECT 124.680 35.100 125.110 37.785 ;
        RECT 125.310 35.985 129.260 37.245 ;
        RECT 129.460 35.100 129.890 37.785 ;
        RECT 134.990 37.445 144.500 37.875 ;
        RECT 134.990 35.040 135.420 37.445 ;
        RECT 135.620 36.010 143.870 37.270 ;
        RECT 144.070 35.040 144.500 37.445 ;
        RECT 64.570 31.890 94.740 32.320 ;
        RECT 64.570 28.470 94.740 28.900 ;
        RECT 64.570 23.890 65.000 28.470 ;
        RECT 65.560 27.170 93.750 27.930 ;
        RECT 65.160 24.430 94.150 25.190 ;
        RECT 94.310 23.890 94.740 28.470 ;
      LAYER nwell ;
        RECT 124.630 25.680 129.940 34.880 ;
        RECT 134.940 27.550 144.550 34.940 ;
      LAYER pwell ;
        RECT 64.570 23.460 94.740 23.890 ;
        RECT 124.680 22.775 125.110 25.460 ;
        RECT 125.310 23.315 129.260 24.575 ;
        RECT 129.460 22.775 129.890 25.460 ;
        RECT 134.990 25.045 135.420 27.450 ;
        RECT 135.620 25.220 143.870 26.480 ;
        RECT 144.070 25.045 144.500 27.450 ;
        RECT 134.990 24.615 144.500 25.045 ;
        RECT 124.680 22.345 129.890 22.775 ;
      LAYER nwell ;
        RECT 69.010 19.010 90.240 22.310 ;
      LAYER pwell ;
        RECT 94.010 20.945 118.580 21.375 ;
        RECT 94.010 18.540 94.440 20.945 ;
        RECT 94.640 19.985 117.950 20.745 ;
        RECT 118.150 18.540 118.580 20.945 ;
      LAYER nwell ;
        RECT 134.940 18.530 144.550 22.490 ;
      LAYER pwell ;
        RECT 55.850 17.575 65.300 18.005 ;
        RECT 55.850 15.735 56.280 17.575 ;
        RECT 56.480 16.275 64.670 17.035 ;
        RECT 64.870 15.735 65.300 17.575 ;
        RECT 55.850 15.305 65.300 15.735 ;
        RECT 69.060 17.575 90.190 18.005 ;
        RECT 69.060 15.735 69.490 17.575 ;
        RECT 69.690 16.275 89.560 17.035 ;
        RECT 89.760 15.735 90.190 17.575 ;
        RECT 69.060 15.305 90.190 15.735 ;
      LAYER nwell ;
        RECT 93.960 14.505 118.630 18.465 ;
      LAYER pwell ;
        RECT 134.990 16.025 135.420 18.430 ;
        RECT 135.620 16.200 143.870 17.460 ;
        RECT 144.070 16.025 144.500 18.430 ;
        RECT 134.990 15.595 144.500 16.025 ;
      LAYER nwell ;
        RECT 93.960 13.890 95.830 14.505 ;
        RECT 55.800 7.000 95.830 13.890 ;
      LAYER li1 ;
        RECT 137.170 77.925 147.200 78.095 ;
        RECT 42.770 76.680 130.840 76.850 ;
        RECT 42.770 73.010 42.940 76.680 ;
        RECT 43.820 76.050 45.430 76.380 ;
        RECT 46.100 76.050 47.710 76.380 ;
        RECT 48.380 76.050 49.990 76.380 ;
        RECT 50.660 76.050 52.270 76.380 ;
        RECT 52.940 76.050 54.550 76.380 ;
        RECT 55.220 76.050 56.830 76.380 ;
        RECT 57.500 76.050 59.110 76.380 ;
        RECT 59.780 76.050 61.390 76.380 ;
        RECT 62.060 76.050 63.670 76.380 ;
        RECT 64.340 76.050 65.950 76.380 ;
        RECT 66.620 76.050 68.230 76.380 ;
        RECT 68.900 76.050 70.510 76.380 ;
        RECT 71.180 76.050 72.790 76.380 ;
        RECT 73.460 76.050 75.070 76.380 ;
        RECT 75.740 76.050 77.350 76.380 ;
        RECT 78.020 76.050 79.630 76.380 ;
        RECT 80.300 76.050 81.910 76.380 ;
        RECT 82.580 76.050 84.190 76.380 ;
        RECT 84.860 76.050 86.470 76.380 ;
        RECT 87.140 76.050 88.750 76.380 ;
        RECT 89.420 76.050 91.030 76.380 ;
        RECT 91.700 76.050 93.310 76.380 ;
        RECT 93.980 76.050 95.590 76.380 ;
        RECT 96.260 76.050 97.870 76.380 ;
        RECT 98.540 76.050 100.150 76.380 ;
        RECT 100.820 76.050 102.430 76.380 ;
        RECT 103.100 76.050 104.710 76.380 ;
        RECT 105.380 76.050 106.990 76.380 ;
        RECT 107.660 76.050 109.270 76.380 ;
        RECT 109.940 76.050 111.550 76.380 ;
        RECT 112.220 76.050 113.830 76.380 ;
        RECT 114.500 76.050 116.110 76.380 ;
        RECT 116.780 76.050 118.390 76.380 ;
        RECT 119.060 76.050 120.670 76.380 ;
        RECT 121.340 76.050 122.950 76.380 ;
        RECT 123.620 76.050 125.230 76.380 ;
        RECT 125.900 76.050 127.510 76.380 ;
        RECT 128.180 76.050 129.790 76.380 ;
        RECT 43.400 75.180 43.570 75.880 ;
        RECT 45.680 75.180 45.850 75.880 ;
        RECT 47.960 75.180 48.130 75.880 ;
        RECT 50.240 75.180 50.410 75.880 ;
        RECT 52.520 75.180 52.690 75.880 ;
        RECT 54.800 75.180 54.970 75.880 ;
        RECT 57.080 75.180 57.250 75.880 ;
        RECT 59.360 75.180 59.530 75.880 ;
        RECT 61.640 75.180 61.810 75.880 ;
        RECT 63.920 75.180 64.090 75.880 ;
        RECT 66.200 75.180 66.370 75.880 ;
        RECT 68.480 75.180 68.650 75.880 ;
        RECT 70.760 75.180 70.930 75.880 ;
        RECT 73.040 75.180 73.210 75.880 ;
        RECT 75.320 75.180 75.490 75.880 ;
        RECT 77.600 75.180 77.770 75.880 ;
        RECT 79.880 75.180 80.050 75.880 ;
        RECT 82.160 75.180 82.330 75.880 ;
        RECT 84.440 75.180 84.610 75.880 ;
        RECT 86.720 75.180 86.890 75.880 ;
        RECT 89.000 75.180 89.170 75.880 ;
        RECT 91.280 75.180 91.450 75.880 ;
        RECT 93.560 75.180 93.730 75.880 ;
        RECT 95.840 75.180 96.010 75.880 ;
        RECT 98.120 75.180 98.290 75.880 ;
        RECT 100.400 75.180 100.570 75.880 ;
        RECT 102.680 75.180 102.850 75.880 ;
        RECT 104.960 75.180 105.130 75.880 ;
        RECT 107.240 75.180 107.410 75.880 ;
        RECT 109.520 75.180 109.690 75.880 ;
        RECT 111.800 75.180 111.970 75.880 ;
        RECT 114.080 75.180 114.250 75.880 ;
        RECT 116.360 75.180 116.530 75.880 ;
        RECT 118.640 75.180 118.810 75.880 ;
        RECT 120.920 75.180 121.090 75.880 ;
        RECT 123.200 75.180 123.370 75.880 ;
        RECT 125.480 75.180 125.650 75.880 ;
        RECT 127.760 75.180 127.930 75.880 ;
        RECT 130.040 75.180 130.210 75.880 ;
        RECT 48.380 74.680 49.990 75.010 ;
        RECT 50.660 74.680 52.270 75.010 ;
        RECT 52.940 74.680 54.550 75.010 ;
        RECT 55.220 74.680 56.830 75.010 ;
        RECT 57.500 74.680 59.110 75.010 ;
        RECT 59.780 74.680 61.390 75.010 ;
        RECT 62.060 74.680 63.670 75.010 ;
        RECT 64.340 74.680 65.950 75.010 ;
        RECT 66.620 74.680 68.230 75.010 ;
        RECT 68.900 74.680 70.510 75.010 ;
        RECT 71.180 74.680 72.790 75.010 ;
        RECT 73.460 74.680 75.070 75.010 ;
        RECT 75.740 74.680 77.350 75.010 ;
        RECT 78.020 74.680 79.630 75.010 ;
        RECT 80.300 74.680 81.910 75.010 ;
        RECT 82.580 74.680 84.190 75.010 ;
        RECT 84.860 74.680 86.470 75.010 ;
        RECT 87.140 74.680 88.750 75.010 ;
        RECT 89.420 74.680 91.030 75.010 ;
        RECT 91.700 74.680 93.310 75.010 ;
        RECT 93.980 74.680 95.590 75.010 ;
        RECT 96.260 74.680 97.870 75.010 ;
        RECT 98.540 74.680 100.150 75.010 ;
        RECT 100.820 74.680 102.430 75.010 ;
        RECT 103.100 74.680 104.710 75.010 ;
        RECT 105.380 74.680 106.990 75.010 ;
        RECT 107.660 74.680 109.270 75.010 ;
        RECT 109.940 74.680 111.550 75.010 ;
        RECT 112.220 74.680 113.830 75.010 ;
        RECT 114.500 74.680 116.110 75.010 ;
        RECT 128.180 74.680 129.790 75.010 ;
        RECT 43.400 73.810 43.570 74.510 ;
        RECT 45.680 73.810 45.850 74.510 ;
        RECT 47.960 73.810 48.130 74.510 ;
        RECT 50.240 73.810 50.410 74.510 ;
        RECT 52.520 73.810 52.690 74.510 ;
        RECT 54.800 73.810 54.970 74.510 ;
        RECT 57.080 73.810 57.250 74.510 ;
        RECT 59.360 73.810 59.530 74.510 ;
        RECT 61.640 73.810 61.810 74.510 ;
        RECT 63.920 73.810 64.090 74.510 ;
        RECT 66.200 73.810 66.370 74.510 ;
        RECT 68.480 73.810 68.650 74.510 ;
        RECT 70.760 73.810 70.930 74.510 ;
        RECT 73.040 73.810 73.210 74.510 ;
        RECT 75.320 73.810 75.490 74.510 ;
        RECT 77.600 73.810 77.770 74.510 ;
        RECT 79.880 73.810 80.050 74.510 ;
        RECT 82.160 73.810 82.330 74.510 ;
        RECT 84.440 73.810 84.610 74.510 ;
        RECT 86.720 73.810 86.890 74.510 ;
        RECT 89.000 73.810 89.170 74.510 ;
        RECT 91.280 73.810 91.450 74.510 ;
        RECT 93.560 73.810 93.730 74.510 ;
        RECT 95.840 73.810 96.010 74.510 ;
        RECT 98.120 73.810 98.290 74.510 ;
        RECT 100.400 73.810 100.570 74.510 ;
        RECT 102.680 73.810 102.850 74.510 ;
        RECT 104.960 73.810 105.130 74.510 ;
        RECT 107.240 73.810 107.410 74.510 ;
        RECT 109.520 73.810 109.690 74.510 ;
        RECT 111.800 73.810 111.970 74.510 ;
        RECT 114.080 73.810 114.250 74.510 ;
        RECT 116.360 73.810 116.530 74.510 ;
        RECT 118.640 73.810 118.810 74.510 ;
        RECT 120.920 73.810 121.090 74.510 ;
        RECT 123.200 73.810 123.370 74.510 ;
        RECT 125.480 73.810 125.650 74.510 ;
        RECT 127.760 73.810 127.930 74.510 ;
        RECT 130.040 73.810 130.210 74.510 ;
        RECT 43.820 73.310 45.430 73.640 ;
        RECT 46.100 73.310 47.710 73.640 ;
        RECT 48.380 73.310 49.990 73.640 ;
        RECT 50.660 73.310 52.270 73.640 ;
        RECT 52.940 73.310 54.550 73.640 ;
        RECT 55.220 73.310 56.830 73.640 ;
        RECT 57.500 73.310 59.110 73.640 ;
        RECT 59.780 73.310 61.390 73.640 ;
        RECT 62.060 73.310 63.670 73.640 ;
        RECT 64.340 73.310 65.950 73.640 ;
        RECT 66.620 73.310 68.230 73.640 ;
        RECT 68.900 73.310 70.510 73.640 ;
        RECT 71.180 73.310 72.790 73.640 ;
        RECT 73.460 73.310 75.070 73.640 ;
        RECT 75.740 73.310 77.350 73.640 ;
        RECT 78.020 73.310 79.630 73.640 ;
        RECT 80.300 73.310 81.910 73.640 ;
        RECT 82.580 73.310 84.190 73.640 ;
        RECT 84.860 73.310 86.470 73.640 ;
        RECT 87.140 73.310 88.750 73.640 ;
        RECT 89.420 73.310 91.030 73.640 ;
        RECT 91.700 73.310 93.310 73.640 ;
        RECT 93.980 73.310 95.590 73.640 ;
        RECT 96.260 73.310 97.870 73.640 ;
        RECT 98.540 73.310 100.150 73.640 ;
        RECT 100.820 73.310 102.430 73.640 ;
        RECT 103.100 73.310 104.710 73.640 ;
        RECT 105.380 73.310 106.990 73.640 ;
        RECT 107.660 73.310 109.270 73.640 ;
        RECT 109.940 73.310 111.550 73.640 ;
        RECT 112.220 73.310 113.830 73.640 ;
        RECT 114.500 73.310 116.110 73.640 ;
        RECT 116.780 73.310 118.390 73.640 ;
        RECT 119.060 73.310 120.670 73.640 ;
        RECT 121.340 73.310 122.950 73.640 ;
        RECT 123.620 73.310 125.230 73.640 ;
        RECT 125.900 73.310 127.510 73.640 ;
        RECT 128.180 73.310 129.790 73.640 ;
        RECT 130.670 73.010 130.840 76.680 ;
        RECT 137.170 75.625 137.340 77.925 ;
        RECT 141.670 77.295 141.840 77.625 ;
        RECT 142.530 77.295 142.700 77.625 ;
        RECT 137.800 76.425 137.970 77.125 ;
        RECT 138.230 76.425 138.400 77.125 ;
        RECT 138.660 76.425 138.830 77.125 ;
        RECT 139.090 76.425 139.260 77.125 ;
        RECT 139.520 76.425 139.690 77.125 ;
        RECT 139.950 76.425 140.120 77.125 ;
        RECT 140.380 76.425 140.550 77.125 ;
        RECT 140.810 76.425 140.980 77.125 ;
        RECT 141.240 76.425 141.410 77.125 ;
        RECT 141.670 76.425 141.840 77.125 ;
        RECT 142.100 76.425 142.270 77.125 ;
        RECT 142.530 76.425 142.700 77.125 ;
        RECT 142.960 76.425 143.130 77.125 ;
        RECT 143.390 76.425 143.560 77.125 ;
        RECT 143.820 76.425 143.990 77.125 ;
        RECT 144.250 76.425 144.420 77.125 ;
        RECT 144.680 76.425 144.850 77.125 ;
        RECT 145.110 76.425 145.280 77.125 ;
        RECT 145.540 76.425 145.710 77.125 ;
        RECT 145.970 76.425 146.140 77.125 ;
        RECT 146.400 76.425 146.570 77.125 ;
        RECT 138.230 75.925 138.400 76.255 ;
        RECT 139.090 75.925 139.260 76.255 ;
        RECT 139.950 75.925 140.120 76.255 ;
        RECT 140.810 75.925 140.980 76.255 ;
        RECT 143.390 75.925 143.560 76.255 ;
        RECT 144.250 75.925 144.420 76.255 ;
        RECT 145.110 75.925 145.280 76.255 ;
        RECT 145.970 75.925 146.140 76.255 ;
        RECT 147.030 75.625 147.200 77.925 ;
        RECT 137.170 75.455 147.200 75.625 ;
        RECT 42.770 72.840 130.840 73.010 ;
        RECT 137.130 74.655 142.080 74.825 ;
        RECT 89.560 71.965 97.870 72.135 ;
        RECT 89.560 69.365 89.730 71.965 ;
        RECT 93.200 71.335 93.370 71.665 ;
        RECT 94.060 71.335 94.230 71.665 ;
        RECT 90.190 70.165 90.360 71.165 ;
        RECT 90.620 70.165 90.790 71.165 ;
        RECT 91.050 70.165 91.220 71.165 ;
        RECT 91.480 70.165 91.650 71.165 ;
        RECT 91.910 70.165 92.080 71.165 ;
        RECT 92.340 70.165 92.510 71.165 ;
        RECT 92.770 70.165 92.940 71.165 ;
        RECT 93.200 70.165 93.370 71.165 ;
        RECT 93.630 70.165 93.800 71.165 ;
        RECT 94.060 70.165 94.230 71.165 ;
        RECT 94.490 70.165 94.660 71.165 ;
        RECT 94.920 70.165 95.090 71.165 ;
        RECT 95.350 70.165 95.520 71.165 ;
        RECT 95.780 70.165 95.950 71.165 ;
        RECT 96.210 70.165 96.380 71.165 ;
        RECT 96.640 70.165 96.810 71.165 ;
        RECT 97.070 70.165 97.240 71.165 ;
        RECT 90.620 69.665 90.790 69.995 ;
        RECT 91.480 69.665 91.650 69.995 ;
        RECT 92.340 69.665 92.510 69.995 ;
        RECT 94.920 69.665 95.090 69.995 ;
        RECT 95.780 69.665 95.950 69.995 ;
        RECT 96.640 69.665 96.810 69.995 ;
        RECT 97.700 69.365 97.870 71.965 ;
        RECT 89.560 69.195 97.870 69.365 ;
        RECT 123.760 71.965 132.070 72.135 ;
        RECT 123.760 69.365 123.930 71.965 ;
        RECT 127.400 71.335 127.570 71.665 ;
        RECT 128.260 71.335 128.430 71.665 ;
        RECT 124.390 70.165 124.560 71.165 ;
        RECT 124.820 70.165 124.990 71.165 ;
        RECT 125.250 70.165 125.420 71.165 ;
        RECT 125.680 70.165 125.850 71.165 ;
        RECT 126.110 70.165 126.280 71.165 ;
        RECT 126.540 70.165 126.710 71.165 ;
        RECT 126.970 70.165 127.140 71.165 ;
        RECT 127.400 70.165 127.570 71.165 ;
        RECT 127.830 70.165 128.000 71.165 ;
        RECT 128.260 70.165 128.430 71.165 ;
        RECT 128.690 70.165 128.860 71.165 ;
        RECT 129.120 70.165 129.290 71.165 ;
        RECT 129.550 70.165 129.720 71.165 ;
        RECT 129.980 70.165 130.150 71.165 ;
        RECT 130.410 70.165 130.580 71.165 ;
        RECT 130.840 70.165 131.010 71.165 ;
        RECT 131.270 70.165 131.440 71.165 ;
        RECT 124.820 69.665 124.990 69.995 ;
        RECT 125.680 69.665 125.850 69.995 ;
        RECT 126.540 69.665 126.710 69.995 ;
        RECT 129.120 69.665 129.290 69.995 ;
        RECT 129.980 69.665 130.150 69.995 ;
        RECT 130.840 69.665 131.010 69.995 ;
        RECT 131.900 69.365 132.070 71.965 ;
        RECT 137.130 69.640 137.300 74.655 ;
        RECT 139.090 74.025 139.260 74.355 ;
        RECT 139.950 74.025 140.120 74.355 ;
        RECT 137.800 73.155 137.970 73.855 ;
        RECT 138.230 73.155 138.400 73.855 ;
        RECT 138.660 73.155 138.830 73.855 ;
        RECT 139.090 73.155 139.260 73.855 ;
        RECT 139.520 73.155 139.690 73.855 ;
        RECT 139.950 73.155 140.120 73.855 ;
        RECT 140.380 73.155 140.550 73.855 ;
        RECT 140.810 73.155 140.980 73.855 ;
        RECT 141.240 73.155 141.410 73.855 ;
        RECT 138.230 72.655 138.400 72.985 ;
        RECT 140.810 72.655 140.980 72.985 ;
        RECT 139.090 71.310 139.260 71.640 ;
        RECT 139.950 71.310 140.120 71.640 ;
        RECT 137.800 70.440 137.970 71.140 ;
        RECT 138.230 70.440 138.400 71.140 ;
        RECT 138.660 70.440 138.830 71.140 ;
        RECT 139.090 70.440 139.260 71.140 ;
        RECT 139.520 70.440 139.690 71.140 ;
        RECT 139.950 70.440 140.120 71.140 ;
        RECT 140.380 70.440 140.550 71.140 ;
        RECT 140.810 70.440 140.980 71.140 ;
        RECT 141.240 70.440 141.410 71.140 ;
        RECT 138.230 69.940 138.400 70.270 ;
        RECT 140.810 69.940 140.980 70.270 ;
        RECT 141.910 69.640 142.080 74.655 ;
        RECT 137.130 69.470 142.080 69.640 ;
        RECT 142.420 74.655 147.290 74.825 ;
        RECT 142.420 69.640 142.590 74.655 ;
        RECT 144.340 74.025 144.510 74.355 ;
        RECT 145.200 74.025 145.370 74.355 ;
        RECT 143.050 73.155 143.220 73.855 ;
        RECT 143.480 73.155 143.650 73.855 ;
        RECT 143.910 73.155 144.080 73.855 ;
        RECT 144.340 73.155 144.510 73.855 ;
        RECT 144.770 73.155 144.940 73.855 ;
        RECT 145.200 73.155 145.370 73.855 ;
        RECT 145.630 73.155 145.800 73.855 ;
        RECT 146.060 73.155 146.230 73.855 ;
        RECT 146.490 73.155 146.660 73.855 ;
        RECT 143.480 72.655 143.650 72.985 ;
        RECT 146.060 72.655 146.230 72.985 ;
        RECT 144.340 71.310 144.510 71.640 ;
        RECT 145.200 71.310 145.370 71.640 ;
        RECT 143.050 70.440 143.220 71.140 ;
        RECT 143.480 70.440 143.650 71.140 ;
        RECT 143.910 70.440 144.080 71.140 ;
        RECT 144.340 70.440 144.510 71.140 ;
        RECT 144.770 70.440 144.940 71.140 ;
        RECT 145.200 70.440 145.370 71.140 ;
        RECT 145.630 70.440 145.800 71.140 ;
        RECT 146.060 70.440 146.230 71.140 ;
        RECT 146.490 70.440 146.660 71.140 ;
        RECT 143.480 69.940 143.650 70.270 ;
        RECT 146.060 69.940 146.230 70.270 ;
        RECT 147.120 69.640 147.290 74.655 ;
        RECT 142.420 69.470 147.290 69.640 ;
        RECT 123.760 69.195 132.070 69.365 ;
        RECT 89.325 68.395 93.335 68.565 ;
        RECT 89.325 66.095 89.495 68.395 ;
        RECT 90.385 67.765 90.555 68.095 ;
        RECT 92.105 67.765 92.275 68.095 ;
        RECT 89.955 66.895 90.125 67.595 ;
        RECT 90.385 66.895 90.555 67.595 ;
        RECT 90.815 66.895 90.985 67.595 ;
        RECT 91.245 66.895 91.415 67.595 ;
        RECT 91.675 66.895 91.845 67.595 ;
        RECT 92.105 66.895 92.275 67.595 ;
        RECT 92.535 66.895 92.705 67.595 ;
        RECT 91.245 66.395 91.415 66.725 ;
        RECT 93.165 66.095 93.335 68.395 ;
        RECT 89.325 65.925 93.335 66.095 ;
        RECT 93.955 68.395 98.045 68.565 ;
        RECT 93.955 66.095 94.125 68.395 ;
        RECT 95.915 67.765 96.085 68.095 ;
        RECT 94.625 66.895 94.795 67.595 ;
        RECT 95.055 66.895 95.225 67.595 ;
        RECT 95.485 66.895 95.655 67.595 ;
        RECT 95.915 66.895 96.085 67.595 ;
        RECT 96.345 66.895 96.515 67.595 ;
        RECT 96.775 66.895 96.945 67.595 ;
        RECT 97.205 66.895 97.375 67.595 ;
        RECT 95.055 66.395 95.225 66.725 ;
        RECT 96.775 66.395 96.945 66.725 ;
        RECT 97.875 66.095 98.045 68.395 ;
        RECT 93.955 65.925 98.045 66.095 ;
        RECT 123.525 68.395 127.535 68.565 ;
        RECT 123.525 66.095 123.695 68.395 ;
        RECT 124.585 67.765 124.755 68.095 ;
        RECT 126.305 67.765 126.475 68.095 ;
        RECT 124.155 66.895 124.325 67.595 ;
        RECT 124.585 66.895 124.755 67.595 ;
        RECT 125.015 66.895 125.185 67.595 ;
        RECT 125.445 66.895 125.615 67.595 ;
        RECT 125.875 66.895 126.045 67.595 ;
        RECT 126.305 66.895 126.475 67.595 ;
        RECT 126.735 66.895 126.905 67.595 ;
        RECT 125.445 66.395 125.615 66.725 ;
        RECT 127.365 66.095 127.535 68.395 ;
        RECT 123.525 65.925 127.535 66.095 ;
        RECT 128.155 68.395 132.245 68.565 ;
        RECT 128.155 66.095 128.325 68.395 ;
        RECT 130.115 67.765 130.285 68.095 ;
        RECT 128.825 66.895 128.995 67.595 ;
        RECT 129.255 66.895 129.425 67.595 ;
        RECT 129.685 66.895 129.855 67.595 ;
        RECT 130.115 66.895 130.285 67.595 ;
        RECT 130.545 66.895 130.715 67.595 ;
        RECT 130.975 66.895 131.145 67.595 ;
        RECT 131.405 66.895 131.575 67.595 ;
        RECT 129.255 66.395 129.425 66.725 ;
        RECT 130.975 66.395 131.145 66.725 ;
        RECT 132.075 66.095 132.245 68.395 ;
        RECT 128.155 65.925 132.245 66.095 ;
        RECT 136.850 68.245 147.480 68.415 ;
        RECT 136.850 65.945 137.020 68.245 ;
        RECT 137.940 67.615 139.550 67.945 ;
        RECT 144.780 67.615 146.390 67.945 ;
        RECT 137.520 66.745 137.690 67.445 ;
        RECT 139.800 66.745 139.970 67.445 ;
        RECT 142.080 66.745 142.250 67.445 ;
        RECT 144.360 66.745 144.530 67.445 ;
        RECT 146.640 66.745 146.810 67.445 ;
        RECT 140.220 66.245 141.830 66.575 ;
        RECT 142.500 66.245 144.110 66.575 ;
        RECT 147.310 65.945 147.480 68.245 ;
        RECT 136.850 65.775 147.480 65.945 ;
        RECT 33.580 65.005 38.530 65.175 ;
        RECT 33.580 61.575 33.750 65.005 ;
        RECT 34.250 62.545 34.420 64.545 ;
        RECT 34.680 62.545 34.850 64.545 ;
        RECT 35.110 62.545 35.280 64.545 ;
        RECT 35.540 62.545 35.710 64.545 ;
        RECT 35.970 62.545 36.140 64.545 ;
        RECT 36.400 62.545 36.570 64.545 ;
        RECT 36.830 62.545 37.000 64.545 ;
        RECT 37.260 62.545 37.430 64.545 ;
        RECT 37.690 62.545 37.860 64.545 ;
        RECT 34.500 62.045 35.030 62.375 ;
        RECT 35.360 62.045 35.890 62.375 ;
        RECT 36.220 62.045 36.750 62.375 ;
        RECT 37.080 62.045 37.610 62.375 ;
        RECT 38.360 61.575 38.530 65.005 ;
        RECT 42.730 64.845 144.560 65.015 ;
        RECT 33.580 58.760 33.750 61.165 ;
        RECT 34.500 60.365 35.030 60.695 ;
        RECT 35.360 60.365 35.890 60.695 ;
        RECT 36.220 60.365 36.750 60.695 ;
        RECT 37.080 60.365 37.610 60.695 ;
        RECT 34.250 59.195 34.420 60.195 ;
        RECT 34.680 59.195 34.850 60.195 ;
        RECT 35.110 59.195 35.280 60.195 ;
        RECT 35.540 59.195 35.710 60.195 ;
        RECT 35.970 59.195 36.140 60.195 ;
        RECT 36.400 59.195 36.570 60.195 ;
        RECT 36.830 59.195 37.000 60.195 ;
        RECT 37.260 59.195 37.430 60.195 ;
        RECT 37.690 59.195 37.860 60.195 ;
        RECT 38.360 58.760 38.530 61.165 ;
        RECT 42.730 59.805 42.900 64.845 ;
        RECT 43.400 63.345 43.570 64.045 ;
        RECT 45.680 63.345 45.850 64.045 ;
        RECT 47.960 63.345 48.130 64.045 ;
        RECT 50.240 63.345 50.410 64.045 ;
        RECT 52.520 63.345 52.690 64.045 ;
        RECT 54.800 63.345 54.970 64.045 ;
        RECT 57.080 63.345 57.250 64.045 ;
        RECT 59.360 63.345 59.530 64.045 ;
        RECT 61.640 63.345 61.810 64.045 ;
        RECT 63.920 63.345 64.090 64.045 ;
        RECT 66.200 63.345 66.370 64.045 ;
        RECT 68.480 63.345 68.650 64.045 ;
        RECT 70.760 63.345 70.930 64.045 ;
        RECT 73.040 63.345 73.210 64.045 ;
        RECT 75.320 63.345 75.490 64.045 ;
        RECT 77.600 63.345 77.770 64.045 ;
        RECT 79.880 63.345 80.050 64.045 ;
        RECT 82.160 63.345 82.330 64.045 ;
        RECT 84.440 63.345 84.610 64.045 ;
        RECT 86.720 63.345 86.890 64.045 ;
        RECT 89.000 63.345 89.170 64.045 ;
        RECT 91.280 63.345 91.450 64.045 ;
        RECT 93.560 63.345 93.730 64.045 ;
        RECT 95.840 63.345 96.010 64.045 ;
        RECT 98.120 63.345 98.290 64.045 ;
        RECT 100.400 63.345 100.570 64.045 ;
        RECT 102.680 63.345 102.850 64.045 ;
        RECT 104.960 63.345 105.130 64.045 ;
        RECT 107.240 63.345 107.410 64.045 ;
        RECT 109.520 63.345 109.690 64.045 ;
        RECT 111.800 63.345 111.970 64.045 ;
        RECT 114.080 63.345 114.250 64.045 ;
        RECT 116.360 63.345 116.530 64.045 ;
        RECT 118.640 63.345 118.810 64.045 ;
        RECT 120.920 63.345 121.090 64.045 ;
        RECT 123.200 63.345 123.370 64.045 ;
        RECT 125.480 63.345 125.650 64.045 ;
        RECT 127.760 63.345 127.930 64.045 ;
        RECT 130.040 63.345 130.210 64.045 ;
        RECT 132.320 63.345 132.490 64.045 ;
        RECT 134.600 63.345 134.770 64.045 ;
        RECT 136.880 63.345 137.050 64.045 ;
        RECT 139.160 63.345 139.330 64.045 ;
        RECT 141.440 63.345 141.610 64.045 ;
        RECT 143.720 63.345 143.890 64.045 ;
        RECT 43.820 62.845 45.430 63.175 ;
        RECT 46.100 62.845 47.710 63.175 ;
        RECT 48.380 62.845 49.990 63.175 ;
        RECT 50.660 62.845 52.270 63.175 ;
        RECT 52.940 62.845 54.550 63.175 ;
        RECT 55.220 62.845 56.830 63.175 ;
        RECT 57.500 62.845 59.110 63.175 ;
        RECT 59.780 62.845 61.390 63.175 ;
        RECT 62.060 62.845 63.670 63.175 ;
        RECT 64.340 62.845 65.950 63.175 ;
        RECT 66.620 62.845 68.230 63.175 ;
        RECT 68.900 62.845 70.510 63.175 ;
        RECT 71.180 62.845 72.790 63.175 ;
        RECT 73.460 62.845 75.070 63.175 ;
        RECT 75.740 62.845 77.350 63.175 ;
        RECT 78.020 62.845 79.630 63.175 ;
        RECT 80.300 62.845 81.910 63.175 ;
        RECT 82.580 62.845 84.190 63.175 ;
        RECT 84.860 62.845 86.470 63.175 ;
        RECT 87.140 62.845 88.750 63.175 ;
        RECT 89.420 62.845 91.030 63.175 ;
        RECT 91.700 62.845 93.310 63.175 ;
        RECT 93.980 62.845 95.590 63.175 ;
        RECT 96.260 62.845 97.870 63.175 ;
        RECT 98.540 62.845 100.150 63.175 ;
        RECT 100.820 62.845 102.430 63.175 ;
        RECT 103.100 62.845 104.710 63.175 ;
        RECT 105.380 62.845 106.990 63.175 ;
        RECT 107.660 62.845 109.270 63.175 ;
        RECT 109.940 62.845 111.550 63.175 ;
        RECT 112.220 62.845 113.830 63.175 ;
        RECT 114.500 62.845 116.110 63.175 ;
        RECT 116.780 62.845 118.390 63.175 ;
        RECT 119.060 62.845 120.670 63.175 ;
        RECT 121.340 62.845 122.950 63.175 ;
        RECT 123.620 62.845 125.230 63.175 ;
        RECT 125.900 62.845 127.510 63.175 ;
        RECT 128.180 62.845 129.790 63.175 ;
        RECT 130.460 62.845 132.070 63.175 ;
        RECT 132.740 62.845 134.350 63.175 ;
        RECT 135.020 62.845 136.630 63.175 ;
        RECT 137.300 62.845 138.910 63.175 ;
        RECT 139.580 62.845 141.190 63.175 ;
        RECT 141.860 62.845 143.470 63.175 ;
        RECT 43.400 61.975 43.570 62.675 ;
        RECT 45.680 61.975 45.850 62.675 ;
        RECT 47.960 61.975 48.130 62.675 ;
        RECT 50.240 61.975 50.410 62.675 ;
        RECT 52.520 61.975 52.690 62.675 ;
        RECT 54.800 61.975 54.970 62.675 ;
        RECT 57.080 61.975 57.250 62.675 ;
        RECT 59.360 61.975 59.530 62.675 ;
        RECT 61.640 61.975 61.810 62.675 ;
        RECT 63.920 61.975 64.090 62.675 ;
        RECT 66.200 61.975 66.370 62.675 ;
        RECT 68.480 61.975 68.650 62.675 ;
        RECT 70.760 61.975 70.930 62.675 ;
        RECT 73.040 61.975 73.210 62.675 ;
        RECT 75.320 61.975 75.490 62.675 ;
        RECT 77.600 61.975 77.770 62.675 ;
        RECT 79.880 61.975 80.050 62.675 ;
        RECT 82.160 61.975 82.330 62.675 ;
        RECT 84.440 61.975 84.610 62.675 ;
        RECT 86.720 61.975 86.890 62.675 ;
        RECT 89.000 61.975 89.170 62.675 ;
        RECT 91.280 61.975 91.450 62.675 ;
        RECT 93.560 61.975 93.730 62.675 ;
        RECT 95.840 61.975 96.010 62.675 ;
        RECT 98.120 61.975 98.290 62.675 ;
        RECT 100.400 61.975 100.570 62.675 ;
        RECT 102.680 61.975 102.850 62.675 ;
        RECT 104.960 61.975 105.130 62.675 ;
        RECT 107.240 61.975 107.410 62.675 ;
        RECT 109.520 61.975 109.690 62.675 ;
        RECT 111.800 61.975 111.970 62.675 ;
        RECT 114.080 61.975 114.250 62.675 ;
        RECT 116.360 61.975 116.530 62.675 ;
        RECT 118.640 61.975 118.810 62.675 ;
        RECT 120.920 61.975 121.090 62.675 ;
        RECT 123.200 61.975 123.370 62.675 ;
        RECT 125.480 61.975 125.650 62.675 ;
        RECT 127.760 61.975 127.930 62.675 ;
        RECT 130.040 61.975 130.210 62.675 ;
        RECT 132.320 61.975 132.490 62.675 ;
        RECT 134.600 61.975 134.770 62.675 ;
        RECT 136.880 61.975 137.050 62.675 ;
        RECT 139.160 61.975 139.330 62.675 ;
        RECT 141.440 61.975 141.610 62.675 ;
        RECT 143.720 61.975 143.890 62.675 ;
        RECT 43.820 61.475 45.430 61.805 ;
        RECT 46.100 61.475 47.710 61.805 ;
        RECT 48.380 61.475 49.990 61.805 ;
        RECT 50.660 61.475 52.270 61.805 ;
        RECT 52.940 61.475 54.550 61.805 ;
        RECT 55.220 61.475 56.830 61.805 ;
        RECT 57.500 61.475 59.110 61.805 ;
        RECT 59.780 61.475 61.390 61.805 ;
        RECT 62.060 61.475 63.670 61.805 ;
        RECT 64.340 61.475 65.950 61.805 ;
        RECT 66.620 61.475 68.230 61.805 ;
        RECT 68.900 61.475 70.510 61.805 ;
        RECT 71.180 61.475 72.790 61.805 ;
        RECT 73.460 61.475 75.070 61.805 ;
        RECT 75.740 61.475 77.350 61.805 ;
        RECT 78.020 61.475 79.630 61.805 ;
        RECT 80.300 61.475 81.910 61.805 ;
        RECT 82.580 61.475 84.190 61.805 ;
        RECT 84.860 61.475 86.470 61.805 ;
        RECT 87.140 61.475 88.750 61.805 ;
        RECT 89.420 61.475 91.030 61.805 ;
        RECT 91.700 61.475 93.310 61.805 ;
        RECT 93.980 61.475 95.590 61.805 ;
        RECT 96.260 61.475 97.870 61.805 ;
        RECT 98.540 61.475 100.150 61.805 ;
        RECT 100.820 61.475 102.430 61.805 ;
        RECT 103.100 61.475 104.710 61.805 ;
        RECT 105.380 61.475 106.990 61.805 ;
        RECT 107.660 61.475 109.270 61.805 ;
        RECT 109.940 61.475 111.550 61.805 ;
        RECT 112.220 61.475 113.830 61.805 ;
        RECT 114.500 61.475 116.110 61.805 ;
        RECT 116.780 61.475 118.390 61.805 ;
        RECT 119.060 61.475 120.670 61.805 ;
        RECT 121.340 61.475 122.950 61.805 ;
        RECT 123.620 61.475 125.230 61.805 ;
        RECT 125.900 61.475 127.510 61.805 ;
        RECT 128.180 61.475 129.790 61.805 ;
        RECT 130.460 61.475 132.070 61.805 ;
        RECT 132.740 61.475 134.350 61.805 ;
        RECT 135.020 61.475 136.630 61.805 ;
        RECT 137.300 61.475 138.910 61.805 ;
        RECT 139.580 61.475 141.190 61.805 ;
        RECT 141.860 61.475 143.470 61.805 ;
        RECT 43.400 60.605 43.570 61.305 ;
        RECT 45.680 60.605 45.850 61.305 ;
        RECT 47.960 60.605 48.130 61.305 ;
        RECT 50.240 60.605 50.410 61.305 ;
        RECT 52.520 60.605 52.690 61.305 ;
        RECT 54.800 60.605 54.970 61.305 ;
        RECT 57.080 60.605 57.250 61.305 ;
        RECT 59.360 60.605 59.530 61.305 ;
        RECT 61.640 60.605 61.810 61.305 ;
        RECT 63.920 60.605 64.090 61.305 ;
        RECT 66.200 60.605 66.370 61.305 ;
        RECT 68.480 60.605 68.650 61.305 ;
        RECT 70.760 60.605 70.930 61.305 ;
        RECT 73.040 60.605 73.210 61.305 ;
        RECT 75.320 60.605 75.490 61.305 ;
        RECT 77.600 60.605 77.770 61.305 ;
        RECT 79.880 60.605 80.050 61.305 ;
        RECT 82.160 60.605 82.330 61.305 ;
        RECT 84.440 60.605 84.610 61.305 ;
        RECT 86.720 60.605 86.890 61.305 ;
        RECT 89.000 60.605 89.170 61.305 ;
        RECT 91.280 60.605 91.450 61.305 ;
        RECT 93.560 60.605 93.730 61.305 ;
        RECT 95.840 60.605 96.010 61.305 ;
        RECT 98.120 60.605 98.290 61.305 ;
        RECT 100.400 60.605 100.570 61.305 ;
        RECT 102.680 60.605 102.850 61.305 ;
        RECT 104.960 60.605 105.130 61.305 ;
        RECT 107.240 60.605 107.410 61.305 ;
        RECT 109.520 60.605 109.690 61.305 ;
        RECT 111.800 60.605 111.970 61.305 ;
        RECT 114.080 60.605 114.250 61.305 ;
        RECT 116.360 60.605 116.530 61.305 ;
        RECT 118.640 60.605 118.810 61.305 ;
        RECT 120.920 60.605 121.090 61.305 ;
        RECT 123.200 60.605 123.370 61.305 ;
        RECT 125.480 60.605 125.650 61.305 ;
        RECT 127.760 60.605 127.930 61.305 ;
        RECT 130.040 60.605 130.210 61.305 ;
        RECT 132.320 60.605 132.490 61.305 ;
        RECT 134.600 60.605 134.770 61.305 ;
        RECT 136.880 60.605 137.050 61.305 ;
        RECT 139.160 60.605 139.330 61.305 ;
        RECT 141.440 60.605 141.610 61.305 ;
        RECT 143.720 60.605 143.890 61.305 ;
        RECT 144.390 59.805 144.560 64.845 ;
        RECT 42.730 59.635 144.560 59.805 ;
        RECT 33.580 58.590 38.530 58.760 ;
        RECT 55.980 53.440 95.650 53.610 ;
        RECT 55.980 47.250 56.150 53.440 ;
        RECT 77.710 52.810 79.320 53.140 ;
        RECT 79.990 52.810 81.600 53.140 ;
        RECT 65.890 51.640 66.060 52.640 ;
        RECT 68.170 51.640 68.340 52.640 ;
        RECT 70.450 51.640 70.620 52.640 ;
        RECT 72.730 51.640 72.900 52.640 ;
        RECT 75.010 51.640 75.180 52.640 ;
        RECT 77.290 51.640 77.460 52.640 ;
        RECT 79.570 51.640 79.740 52.640 ;
        RECT 81.850 51.640 82.020 52.640 ;
        RECT 84.130 51.640 84.300 52.640 ;
        RECT 86.410 51.640 86.580 52.640 ;
        RECT 88.690 51.640 88.860 52.640 ;
        RECT 90.970 51.640 91.140 52.640 ;
        RECT 93.250 51.640 93.420 52.640 ;
        RECT 66.310 51.140 67.920 51.470 ;
        RECT 68.590 51.140 70.200 51.470 ;
        RECT 70.870 51.140 72.480 51.470 ;
        RECT 73.150 51.140 74.760 51.470 ;
        RECT 75.430 51.140 77.040 51.470 ;
        RECT 82.270 51.140 83.880 51.470 ;
        RECT 84.550 51.140 86.160 51.470 ;
        RECT 86.830 51.140 88.440 51.470 ;
        RECT 89.110 51.140 90.720 51.470 ;
        RECT 91.390 51.140 93.000 51.470 ;
        RECT 57.070 49.220 57.960 49.550 ;
        RECT 63.190 49.220 64.080 49.550 ;
        RECT 64.750 49.220 65.640 49.550 ;
        RECT 66.310 49.220 67.920 49.550 ;
        RECT 68.590 49.220 70.200 49.550 ;
        RECT 70.870 49.220 72.480 49.550 ;
        RECT 73.150 49.220 74.760 49.550 ;
        RECT 75.430 49.220 77.040 49.550 ;
        RECT 77.710 49.220 79.320 49.550 ;
        RECT 79.990 49.220 81.600 49.550 ;
        RECT 82.270 49.220 83.880 49.550 ;
        RECT 84.550 49.220 86.160 49.550 ;
        RECT 86.830 49.220 88.440 49.550 ;
        RECT 89.110 49.220 90.720 49.550 ;
        RECT 91.390 49.220 93.000 49.550 ;
        RECT 93.670 49.220 94.560 49.550 ;
        RECT 56.650 48.050 56.820 49.050 ;
        RECT 57.430 48.050 57.600 49.050 ;
        RECT 58.210 48.050 58.380 49.050 ;
        RECT 60.490 48.050 60.660 49.050 ;
        RECT 62.770 48.050 62.940 49.050 ;
        RECT 63.550 48.050 63.720 49.050 ;
        RECT 64.330 48.050 64.500 49.050 ;
        RECT 65.110 48.050 65.280 49.050 ;
        RECT 65.890 48.050 66.060 49.050 ;
        RECT 68.170 48.050 68.340 49.050 ;
        RECT 70.450 48.050 70.620 49.050 ;
        RECT 72.730 48.050 72.900 49.050 ;
        RECT 75.010 48.050 75.180 49.050 ;
        RECT 77.290 48.050 77.460 49.050 ;
        RECT 79.570 48.050 79.740 49.050 ;
        RECT 81.850 48.050 82.020 49.050 ;
        RECT 84.130 48.050 84.300 49.050 ;
        RECT 86.410 48.050 86.580 49.050 ;
        RECT 88.690 48.050 88.860 49.050 ;
        RECT 90.970 48.050 91.140 49.050 ;
        RECT 93.250 48.050 93.420 49.050 ;
        RECT 94.030 48.050 94.200 49.050 ;
        RECT 94.810 48.050 94.980 49.050 ;
        RECT 58.630 47.550 60.240 47.880 ;
        RECT 60.910 47.550 62.520 47.880 ;
        RECT 66.310 47.550 67.920 47.880 ;
        RECT 68.590 47.550 70.200 47.880 ;
        RECT 70.870 47.550 72.480 47.880 ;
        RECT 73.150 47.550 74.760 47.880 ;
        RECT 75.430 47.550 77.040 47.880 ;
        RECT 77.710 47.550 79.320 47.880 ;
        RECT 79.990 47.550 81.600 47.880 ;
        RECT 82.270 47.550 83.880 47.880 ;
        RECT 84.550 47.550 86.160 47.880 ;
        RECT 86.830 47.550 88.440 47.880 ;
        RECT 89.110 47.550 90.720 47.880 ;
        RECT 91.390 47.550 93.000 47.880 ;
        RECT 95.480 47.250 95.650 53.440 ;
        RECT 55.980 47.080 95.650 47.250 ;
        RECT 94.140 45.935 118.450 46.105 ;
        RECT 55.980 45.185 65.170 45.355 ;
        RECT 55.980 43.085 56.150 45.185 ;
        RECT 58.630 44.555 60.240 44.885 ;
        RECT 60.910 44.555 62.520 44.885 ;
        RECT 56.650 43.885 56.820 44.385 ;
        RECT 57.430 43.885 57.600 44.385 ;
        RECT 58.210 43.885 58.380 44.385 ;
        RECT 60.490 43.885 60.660 44.385 ;
        RECT 62.770 43.885 62.940 44.385 ;
        RECT 63.550 43.885 63.720 44.385 ;
        RECT 64.330 43.885 64.500 44.385 ;
        RECT 57.070 43.385 57.960 43.715 ;
        RECT 63.190 43.385 64.080 43.715 ;
        RECT 65.000 43.085 65.170 45.185 ;
        RECT 55.980 42.915 65.170 43.085 ;
        RECT 69.190 45.185 90.060 45.355 ;
        RECT 69.190 43.085 69.360 45.185 ;
        RECT 70.245 44.555 72.215 44.885 ;
        RECT 72.840 44.555 74.450 44.885 ;
        RECT 75.120 44.555 76.730 44.885 ;
        RECT 77.365 44.555 79.335 44.885 ;
        RECT 79.925 44.555 81.895 44.885 ;
        RECT 82.520 44.555 84.130 44.885 ;
        RECT 84.800 44.555 86.410 44.885 ;
        RECT 87.045 44.555 89.015 44.885 ;
        RECT 69.860 43.885 70.030 44.385 ;
        RECT 71.140 43.885 71.310 44.385 ;
        RECT 72.420 43.885 72.590 44.385 ;
        RECT 74.700 43.885 74.870 44.385 ;
        RECT 76.980 43.885 77.150 44.385 ;
        RECT 78.260 43.885 78.430 44.385 ;
        RECT 79.540 43.885 79.710 44.385 ;
        RECT 80.820 43.885 80.990 44.385 ;
        RECT 82.100 43.885 82.270 44.385 ;
        RECT 84.380 43.885 84.550 44.385 ;
        RECT 86.660 43.885 86.830 44.385 ;
        RECT 87.940 43.885 88.110 44.385 ;
        RECT 89.220 43.885 89.390 44.385 ;
        RECT 70.245 43.385 72.215 43.715 ;
        RECT 72.840 43.385 74.450 43.715 ;
        RECT 75.120 43.385 76.730 43.715 ;
        RECT 77.365 43.385 79.335 43.715 ;
        RECT 79.925 43.385 81.895 43.715 ;
        RECT 87.045 43.385 89.015 43.715 ;
        RECT 89.890 43.085 90.060 45.185 ;
        RECT 69.190 42.915 90.060 43.085 ;
        RECT 94.140 42.505 94.310 45.935 ;
        RECT 94.810 44.475 94.980 45.475 ;
        RECT 97.090 44.475 97.260 45.475 ;
        RECT 99.370 44.475 99.540 45.475 ;
        RECT 101.650 44.475 101.820 45.475 ;
        RECT 103.930 44.475 104.100 45.475 ;
        RECT 106.210 44.475 106.380 45.475 ;
        RECT 108.490 44.475 108.660 45.475 ;
        RECT 110.770 44.475 110.940 45.475 ;
        RECT 113.050 44.475 113.220 45.475 ;
        RECT 115.330 44.475 115.500 45.475 ;
        RECT 117.610 44.475 117.780 45.475 ;
        RECT 95.230 43.975 96.840 44.305 ;
        RECT 97.510 43.975 99.120 44.305 ;
        RECT 99.790 43.975 101.400 44.305 ;
        RECT 102.070 43.975 103.680 44.305 ;
        RECT 104.350 43.975 105.960 44.305 ;
        RECT 106.630 43.975 108.240 44.305 ;
        RECT 108.910 43.975 110.520 44.305 ;
        RECT 111.190 43.975 112.800 44.305 ;
        RECT 113.470 43.975 115.080 44.305 ;
        RECT 115.750 43.975 117.360 44.305 ;
        RECT 118.280 42.505 118.450 45.935 ;
        RECT 124.460 45.920 129.410 46.090 ;
        RECT 124.460 42.490 124.630 45.920 ;
        RECT 125.130 43.460 125.300 45.460 ;
        RECT 125.560 43.460 125.730 45.460 ;
        RECT 125.990 43.460 126.160 45.460 ;
        RECT 126.420 43.460 126.590 45.460 ;
        RECT 126.850 43.460 127.020 45.460 ;
        RECT 127.280 43.460 127.450 45.460 ;
        RECT 127.710 43.460 127.880 45.460 ;
        RECT 128.140 43.460 128.310 45.460 ;
        RECT 128.570 43.460 128.740 45.460 ;
        RECT 125.380 42.960 125.910 43.290 ;
        RECT 126.240 42.960 126.770 43.290 ;
        RECT 127.100 42.960 127.630 43.290 ;
        RECT 127.960 42.960 128.490 43.290 ;
        RECT 129.240 42.490 129.410 45.920 ;
        RECT 135.120 45.920 144.370 46.090 ;
        RECT 135.120 42.490 135.290 45.920 ;
        RECT 135.790 43.460 135.960 45.460 ;
        RECT 136.220 43.460 136.390 45.460 ;
        RECT 136.650 43.460 136.820 45.460 ;
        RECT 137.080 43.460 137.250 45.460 ;
        RECT 137.510 43.460 137.680 45.460 ;
        RECT 137.940 43.460 138.110 45.460 ;
        RECT 138.370 43.460 138.540 45.460 ;
        RECT 138.800 43.460 138.970 45.460 ;
        RECT 139.230 43.460 139.400 45.460 ;
        RECT 139.660 43.460 139.830 45.460 ;
        RECT 140.090 43.460 140.260 45.460 ;
        RECT 140.520 43.460 140.690 45.460 ;
        RECT 140.950 43.460 141.120 45.460 ;
        RECT 141.380 43.460 141.550 45.460 ;
        RECT 141.810 43.460 141.980 45.460 ;
        RECT 142.240 43.460 142.410 45.460 ;
        RECT 142.670 43.460 142.840 45.460 ;
        RECT 143.100 43.460 143.270 45.460 ;
        RECT 143.530 43.460 143.700 45.460 ;
        RECT 136.040 42.960 136.570 43.290 ;
        RECT 136.900 42.960 137.430 43.290 ;
        RECT 137.760 42.960 138.290 43.290 ;
        RECT 138.620 42.960 139.150 43.290 ;
        RECT 139.480 42.960 140.010 43.290 ;
        RECT 140.340 42.960 140.870 43.290 ;
        RECT 141.200 42.960 141.730 43.290 ;
        RECT 142.060 42.960 142.590 43.290 ;
        RECT 142.920 42.960 143.450 43.290 ;
        RECT 144.200 42.490 144.370 45.920 ;
        RECT 69.190 41.430 90.060 41.600 ;
        RECT 69.190 38.830 69.360 41.430 ;
        RECT 70.245 40.800 72.215 41.130 ;
        RECT 72.840 40.800 74.450 41.130 ;
        RECT 75.120 40.800 76.730 41.130 ;
        RECT 77.365 40.800 79.335 41.130 ;
        RECT 79.925 40.800 81.895 41.130 ;
        RECT 87.045 40.800 89.015 41.130 ;
        RECT 69.860 39.630 70.030 40.630 ;
        RECT 71.140 39.630 71.310 40.630 ;
        RECT 72.420 39.630 72.590 40.630 ;
        RECT 74.700 39.630 74.870 40.630 ;
        RECT 76.980 39.630 77.150 40.630 ;
        RECT 78.260 39.630 78.430 40.630 ;
        RECT 79.540 39.630 79.710 40.630 ;
        RECT 80.820 39.630 80.990 40.630 ;
        RECT 82.100 39.630 82.270 40.630 ;
        RECT 84.380 39.630 84.550 40.630 ;
        RECT 86.660 39.630 86.830 40.630 ;
        RECT 87.940 39.630 88.110 40.630 ;
        RECT 89.220 39.630 89.390 40.630 ;
        RECT 70.245 39.130 72.215 39.460 ;
        RECT 72.840 39.130 74.450 39.460 ;
        RECT 75.120 39.130 76.730 39.460 ;
        RECT 77.365 39.130 79.335 39.460 ;
        RECT 79.925 39.130 81.895 39.460 ;
        RECT 82.520 39.130 84.130 39.460 ;
        RECT 84.800 39.130 86.410 39.460 ;
        RECT 87.045 39.130 89.015 39.460 ;
        RECT 89.890 38.830 90.060 41.430 ;
        RECT 94.140 39.715 94.310 42.120 ;
        RECT 95.230 40.845 96.840 41.175 ;
        RECT 97.510 40.845 99.120 41.175 ;
        RECT 99.790 40.845 101.400 41.175 ;
        RECT 102.070 40.845 103.680 41.175 ;
        RECT 104.350 40.845 105.960 41.175 ;
        RECT 106.630 40.845 108.240 41.175 ;
        RECT 108.910 40.845 110.520 41.175 ;
        RECT 111.190 40.845 112.800 41.175 ;
        RECT 113.470 40.845 115.080 41.175 ;
        RECT 115.750 40.845 117.360 41.175 ;
        RECT 94.810 40.175 94.980 40.675 ;
        RECT 97.090 40.175 97.260 40.675 ;
        RECT 99.370 40.175 99.540 40.675 ;
        RECT 101.650 40.175 101.820 40.675 ;
        RECT 103.930 40.175 104.100 40.675 ;
        RECT 106.210 40.175 106.380 40.675 ;
        RECT 108.490 40.175 108.660 40.675 ;
        RECT 110.770 40.175 110.940 40.675 ;
        RECT 113.050 40.175 113.220 40.675 ;
        RECT 115.330 40.175 115.500 40.675 ;
        RECT 117.610 40.175 117.780 40.675 ;
        RECT 118.280 39.715 118.450 42.120 ;
        RECT 94.140 39.545 118.450 39.715 ;
        RECT 124.460 39.675 124.630 42.080 ;
        RECT 125.380 41.280 125.910 41.610 ;
        RECT 126.240 41.280 126.770 41.610 ;
        RECT 127.100 41.280 127.630 41.610 ;
        RECT 127.960 41.280 128.490 41.610 ;
        RECT 125.130 40.110 125.300 41.110 ;
        RECT 125.560 40.110 125.730 41.110 ;
        RECT 125.990 40.110 126.160 41.110 ;
        RECT 126.420 40.110 126.590 41.110 ;
        RECT 126.850 40.110 127.020 41.110 ;
        RECT 127.280 40.110 127.450 41.110 ;
        RECT 127.710 40.110 127.880 41.110 ;
        RECT 128.140 40.110 128.310 41.110 ;
        RECT 128.570 40.110 128.740 41.110 ;
        RECT 129.240 39.675 129.410 42.080 ;
        RECT 124.460 39.505 129.410 39.675 ;
        RECT 135.120 39.675 135.290 42.080 ;
        RECT 136.040 41.280 136.570 41.610 ;
        RECT 136.900 41.280 137.430 41.610 ;
        RECT 137.760 41.280 138.290 41.610 ;
        RECT 138.620 41.280 139.150 41.610 ;
        RECT 139.480 41.280 140.010 41.610 ;
        RECT 140.340 41.280 140.870 41.610 ;
        RECT 141.200 41.280 141.730 41.610 ;
        RECT 142.060 41.280 142.590 41.610 ;
        RECT 142.920 41.280 143.450 41.610 ;
        RECT 135.790 40.110 135.960 41.110 ;
        RECT 136.220 40.110 136.390 41.110 ;
        RECT 136.650 40.110 136.820 41.110 ;
        RECT 137.080 40.110 137.250 41.110 ;
        RECT 137.510 40.110 137.680 41.110 ;
        RECT 137.940 40.110 138.110 41.110 ;
        RECT 138.370 40.110 138.540 41.110 ;
        RECT 138.800 40.110 138.970 41.110 ;
        RECT 139.230 40.110 139.400 41.110 ;
        RECT 139.660 40.110 139.830 41.110 ;
        RECT 140.090 40.110 140.260 41.110 ;
        RECT 140.520 40.110 140.690 41.110 ;
        RECT 140.950 40.110 141.120 41.110 ;
        RECT 141.380 40.110 141.550 41.110 ;
        RECT 141.810 40.110 141.980 41.110 ;
        RECT 142.240 40.110 142.410 41.110 ;
        RECT 142.670 40.110 142.840 41.110 ;
        RECT 143.100 40.110 143.270 41.110 ;
        RECT 143.530 40.110 143.700 41.110 ;
        RECT 144.200 39.675 144.370 42.080 ;
        RECT 135.120 39.505 144.370 39.675 ;
        RECT 69.190 38.660 90.060 38.830 ;
        RECT 124.810 37.915 129.760 38.085 ;
        RECT 64.700 37.030 94.610 37.200 ;
        RECT 64.700 32.190 64.870 37.030 ;
        RECT 68.310 36.400 69.920 36.730 ;
        RECT 70.590 36.400 72.200 36.730 ;
        RECT 72.870 36.400 74.480 36.730 ;
        RECT 75.150 36.400 76.760 36.730 ;
        RECT 77.395 36.400 79.365 36.730 ;
        RECT 79.955 36.400 81.925 36.730 ;
        RECT 82.550 36.400 84.160 36.730 ;
        RECT 84.830 36.400 86.440 36.730 ;
        RECT 87.110 36.400 88.720 36.730 ;
        RECT 89.390 36.400 91.000 36.730 ;
        RECT 65.330 35.730 65.500 36.230 ;
        RECT 66.610 35.730 66.780 36.230 ;
        RECT 67.890 35.730 68.060 36.230 ;
        RECT 70.170 35.730 70.340 36.230 ;
        RECT 72.450 35.730 72.620 36.230 ;
        RECT 74.730 35.730 74.900 36.230 ;
        RECT 77.010 35.730 77.180 36.230 ;
        RECT 78.290 35.730 78.460 36.230 ;
        RECT 79.570 35.730 79.740 36.230 ;
        RECT 80.850 35.730 81.020 36.230 ;
        RECT 82.130 35.730 82.300 36.230 ;
        RECT 84.410 35.730 84.580 36.230 ;
        RECT 86.690 35.730 86.860 36.230 ;
        RECT 88.970 35.730 89.140 36.230 ;
        RECT 91.250 35.730 91.420 36.230 ;
        RECT 92.530 35.730 92.700 36.230 ;
        RECT 93.810 35.730 93.980 36.230 ;
        RECT 65.715 35.230 67.685 35.560 ;
        RECT 68.310 35.230 69.920 35.560 ;
        RECT 70.590 35.230 72.200 35.560 ;
        RECT 72.870 35.230 74.480 35.560 ;
        RECT 75.150 35.230 76.760 35.560 ;
        RECT 77.395 35.230 79.365 35.560 ;
        RECT 79.955 35.230 81.925 35.560 ;
        RECT 82.550 35.230 84.160 35.560 ;
        RECT 84.830 35.230 86.440 35.560 ;
        RECT 87.110 35.230 88.720 35.560 ;
        RECT 89.390 35.230 91.000 35.560 ;
        RECT 91.635 35.230 93.605 35.560 ;
        RECT 66.115 33.660 68.805 33.990 ;
        RECT 69.395 33.660 72.085 33.990 ;
        RECT 87.235 33.660 89.925 33.990 ;
        RECT 90.515 33.660 93.205 33.990 ;
        RECT 65.730 32.990 65.900 33.490 ;
        RECT 69.010 32.990 69.180 33.490 ;
        RECT 72.290 32.990 72.460 33.490 ;
        RECT 79.570 32.990 79.740 33.490 ;
        RECT 86.850 32.990 87.020 33.490 ;
        RECT 90.130 32.990 90.300 33.490 ;
        RECT 93.410 32.990 93.580 33.490 ;
        RECT 66.115 32.490 68.805 32.820 ;
        RECT 69.395 32.490 72.085 32.820 ;
        RECT 72.690 32.490 79.340 32.820 ;
        RECT 79.970 32.490 86.620 32.820 ;
        RECT 87.235 32.490 89.925 32.820 ;
        RECT 90.515 32.490 93.205 32.820 ;
        RECT 94.440 32.190 94.610 37.030 ;
        RECT 124.810 35.230 124.980 37.915 ;
        RECT 125.730 37.285 126.260 37.615 ;
        RECT 126.590 37.285 127.120 37.615 ;
        RECT 127.450 37.285 127.980 37.615 ;
        RECT 128.310 37.285 128.840 37.615 ;
        RECT 125.480 36.115 125.650 37.115 ;
        RECT 125.910 36.115 126.080 37.115 ;
        RECT 126.340 36.115 126.510 37.115 ;
        RECT 126.770 36.115 126.940 37.115 ;
        RECT 127.200 36.115 127.370 37.115 ;
        RECT 127.630 36.115 127.800 37.115 ;
        RECT 128.060 36.115 128.230 37.115 ;
        RECT 128.490 36.115 128.660 37.115 ;
        RECT 128.920 36.115 129.090 37.115 ;
        RECT 125.730 35.615 126.260 35.945 ;
        RECT 126.590 35.615 127.120 35.945 ;
        RECT 127.450 35.615 127.980 35.945 ;
        RECT 128.310 35.615 128.840 35.945 ;
        RECT 129.590 35.230 129.760 37.915 ;
        RECT 135.120 37.575 144.370 37.745 ;
        RECT 135.120 35.170 135.290 37.575 ;
        RECT 135.790 36.140 135.960 37.140 ;
        RECT 136.220 36.140 136.390 37.140 ;
        RECT 136.650 36.140 136.820 37.140 ;
        RECT 137.080 36.140 137.250 37.140 ;
        RECT 137.510 36.140 137.680 37.140 ;
        RECT 137.940 36.140 138.110 37.140 ;
        RECT 138.370 36.140 138.540 37.140 ;
        RECT 138.800 36.140 138.970 37.140 ;
        RECT 139.230 36.140 139.400 37.140 ;
        RECT 139.660 36.140 139.830 37.140 ;
        RECT 140.090 36.140 140.260 37.140 ;
        RECT 140.520 36.140 140.690 37.140 ;
        RECT 140.950 36.140 141.120 37.140 ;
        RECT 141.380 36.140 141.550 37.140 ;
        RECT 141.810 36.140 141.980 37.140 ;
        RECT 142.240 36.140 142.410 37.140 ;
        RECT 142.670 36.140 142.840 37.140 ;
        RECT 143.100 36.140 143.270 37.140 ;
        RECT 143.530 36.140 143.700 37.140 ;
        RECT 136.040 35.640 136.570 35.970 ;
        RECT 136.900 35.640 137.430 35.970 ;
        RECT 137.760 35.640 138.290 35.970 ;
        RECT 138.620 35.640 139.150 35.970 ;
        RECT 139.480 35.640 140.010 35.970 ;
        RECT 140.340 35.640 140.870 35.970 ;
        RECT 141.200 35.640 141.730 35.970 ;
        RECT 142.060 35.640 142.590 35.970 ;
        RECT 142.920 35.640 143.450 35.970 ;
        RECT 144.200 35.170 144.370 37.575 ;
        RECT 64.700 32.020 94.610 32.190 ;
        RECT 124.810 30.365 124.980 34.700 ;
        RECT 125.730 33.985 126.260 34.315 ;
        RECT 126.590 33.985 127.120 34.315 ;
        RECT 127.450 33.985 127.980 34.315 ;
        RECT 128.310 33.985 128.840 34.315 ;
        RECT 125.480 32.815 125.650 33.815 ;
        RECT 125.910 32.815 126.080 33.815 ;
        RECT 126.340 32.815 126.510 33.815 ;
        RECT 126.770 32.815 126.940 33.815 ;
        RECT 127.200 32.815 127.370 33.815 ;
        RECT 127.630 32.815 127.800 33.815 ;
        RECT 128.060 32.815 128.230 33.815 ;
        RECT 128.490 32.815 128.660 33.815 ;
        RECT 128.920 32.815 129.090 33.815 ;
        RECT 125.480 31.165 125.650 32.165 ;
        RECT 125.910 31.165 126.080 32.165 ;
        RECT 126.340 31.165 126.510 32.165 ;
        RECT 126.770 31.165 126.940 32.165 ;
        RECT 127.200 31.165 127.370 32.165 ;
        RECT 127.630 31.165 127.800 32.165 ;
        RECT 128.060 31.165 128.230 32.165 ;
        RECT 128.490 31.165 128.660 32.165 ;
        RECT 128.920 31.165 129.090 32.165 ;
        RECT 125.730 30.665 126.260 30.995 ;
        RECT 126.590 30.665 127.120 30.995 ;
        RECT 127.450 30.665 127.980 30.995 ;
        RECT 128.310 30.665 128.840 30.995 ;
        RECT 129.590 30.365 129.760 34.700 ;
        RECT 124.810 30.195 129.760 30.365 ;
        RECT 64.700 28.600 94.610 28.770 ;
        RECT 64.700 23.760 64.870 28.600 ;
        RECT 66.115 27.970 68.805 28.300 ;
        RECT 69.395 27.970 72.085 28.300 ;
        RECT 72.690 27.970 79.340 28.300 ;
        RECT 79.970 27.970 86.620 28.300 ;
        RECT 87.235 27.970 89.925 28.300 ;
        RECT 90.515 27.970 93.205 28.300 ;
        RECT 65.730 27.300 65.900 27.800 ;
        RECT 69.010 27.300 69.180 27.800 ;
        RECT 72.290 27.300 72.460 27.800 ;
        RECT 79.570 27.300 79.740 27.800 ;
        RECT 86.850 27.300 87.020 27.800 ;
        RECT 90.130 27.300 90.300 27.800 ;
        RECT 93.410 27.300 93.580 27.800 ;
        RECT 66.115 26.800 68.805 27.130 ;
        RECT 69.395 26.800 72.085 27.130 ;
        RECT 87.235 26.800 89.925 27.130 ;
        RECT 90.515 26.800 93.205 27.130 ;
        RECT 65.715 25.230 67.685 25.560 ;
        RECT 68.310 25.230 69.920 25.560 ;
        RECT 70.590 25.230 72.200 25.560 ;
        RECT 72.870 25.230 74.480 25.560 ;
        RECT 75.150 25.230 76.760 25.560 ;
        RECT 77.395 25.230 79.365 25.560 ;
        RECT 79.955 25.230 81.925 25.560 ;
        RECT 82.550 25.230 84.160 25.560 ;
        RECT 84.830 25.230 86.440 25.560 ;
        RECT 87.110 25.230 88.720 25.560 ;
        RECT 89.390 25.230 91.000 25.560 ;
        RECT 91.635 25.230 93.605 25.560 ;
        RECT 65.330 24.560 65.500 25.060 ;
        RECT 66.610 24.560 66.780 25.060 ;
        RECT 67.890 24.560 68.060 25.060 ;
        RECT 70.170 24.560 70.340 25.060 ;
        RECT 72.450 24.560 72.620 25.060 ;
        RECT 74.730 24.560 74.900 25.060 ;
        RECT 77.010 24.560 77.180 25.060 ;
        RECT 78.290 24.560 78.460 25.060 ;
        RECT 79.570 24.560 79.740 25.060 ;
        RECT 80.850 24.560 81.020 25.060 ;
        RECT 82.130 24.560 82.300 25.060 ;
        RECT 84.410 24.560 84.580 25.060 ;
        RECT 86.690 24.560 86.860 25.060 ;
        RECT 88.970 24.560 89.140 25.060 ;
        RECT 91.250 24.560 91.420 25.060 ;
        RECT 92.530 24.560 92.700 25.060 ;
        RECT 93.810 24.560 93.980 25.060 ;
        RECT 68.310 24.060 69.920 24.390 ;
        RECT 70.590 24.060 72.200 24.390 ;
        RECT 72.870 24.060 74.480 24.390 ;
        RECT 75.150 24.060 76.760 24.390 ;
        RECT 77.395 24.060 79.365 24.390 ;
        RECT 79.955 24.060 81.925 24.390 ;
        RECT 82.550 24.060 84.160 24.390 ;
        RECT 84.830 24.060 86.440 24.390 ;
        RECT 87.110 24.060 88.720 24.390 ;
        RECT 89.390 24.060 91.000 24.390 ;
        RECT 94.440 23.760 94.610 28.600 ;
        RECT 124.810 25.860 124.980 30.195 ;
        RECT 125.730 29.565 126.260 29.895 ;
        RECT 126.590 29.565 127.120 29.895 ;
        RECT 127.450 29.565 127.980 29.895 ;
        RECT 128.310 29.565 128.840 29.895 ;
        RECT 125.480 28.395 125.650 29.395 ;
        RECT 125.910 28.395 126.080 29.395 ;
        RECT 126.340 28.395 126.510 29.395 ;
        RECT 126.770 28.395 126.940 29.395 ;
        RECT 127.200 28.395 127.370 29.395 ;
        RECT 127.630 28.395 127.800 29.395 ;
        RECT 128.060 28.395 128.230 29.395 ;
        RECT 128.490 28.395 128.660 29.395 ;
        RECT 128.920 28.395 129.090 29.395 ;
        RECT 125.480 26.745 125.650 27.745 ;
        RECT 125.910 26.745 126.080 27.745 ;
        RECT 126.340 26.745 126.510 27.745 ;
        RECT 126.770 26.745 126.940 27.745 ;
        RECT 127.200 26.745 127.370 27.745 ;
        RECT 127.630 26.745 127.800 27.745 ;
        RECT 128.060 26.745 128.230 27.745 ;
        RECT 128.490 26.745 128.660 27.745 ;
        RECT 128.920 26.745 129.090 27.745 ;
        RECT 125.730 26.245 126.260 26.575 ;
        RECT 126.590 26.245 127.120 26.575 ;
        RECT 127.450 26.245 127.980 26.575 ;
        RECT 128.310 26.245 128.840 26.575 ;
        RECT 129.590 25.860 129.760 30.195 ;
        RECT 135.120 31.330 135.290 34.760 ;
        RECT 136.040 33.960 136.570 34.290 ;
        RECT 136.900 33.960 137.430 34.290 ;
        RECT 137.760 33.960 138.290 34.290 ;
        RECT 138.620 33.960 139.150 34.290 ;
        RECT 139.480 33.960 140.010 34.290 ;
        RECT 140.340 33.960 140.870 34.290 ;
        RECT 141.200 33.960 141.730 34.290 ;
        RECT 142.060 33.960 142.590 34.290 ;
        RECT 142.920 33.960 143.450 34.290 ;
        RECT 135.790 31.790 135.960 33.790 ;
        RECT 136.220 31.790 136.390 33.790 ;
        RECT 136.650 31.790 136.820 33.790 ;
        RECT 137.080 31.790 137.250 33.790 ;
        RECT 137.510 31.790 137.680 33.790 ;
        RECT 137.940 31.790 138.110 33.790 ;
        RECT 138.370 31.790 138.540 33.790 ;
        RECT 138.800 31.790 138.970 33.790 ;
        RECT 139.230 31.790 139.400 33.790 ;
        RECT 139.660 31.790 139.830 33.790 ;
        RECT 140.090 31.790 140.260 33.790 ;
        RECT 140.520 31.790 140.690 33.790 ;
        RECT 140.950 31.790 141.120 33.790 ;
        RECT 141.380 31.790 141.550 33.790 ;
        RECT 141.810 31.790 141.980 33.790 ;
        RECT 142.240 31.790 142.410 33.790 ;
        RECT 142.670 31.790 142.840 33.790 ;
        RECT 143.100 31.790 143.270 33.790 ;
        RECT 143.530 31.790 143.700 33.790 ;
        RECT 144.200 31.330 144.370 34.760 ;
        RECT 135.120 31.160 144.370 31.330 ;
        RECT 135.120 27.730 135.290 31.160 ;
        RECT 135.790 28.700 135.960 30.700 ;
        RECT 136.220 28.700 136.390 30.700 ;
        RECT 136.650 28.700 136.820 30.700 ;
        RECT 137.080 28.700 137.250 30.700 ;
        RECT 137.510 28.700 137.680 30.700 ;
        RECT 137.940 28.700 138.110 30.700 ;
        RECT 138.370 28.700 138.540 30.700 ;
        RECT 138.800 28.700 138.970 30.700 ;
        RECT 139.230 28.700 139.400 30.700 ;
        RECT 139.660 28.700 139.830 30.700 ;
        RECT 140.090 28.700 140.260 30.700 ;
        RECT 140.520 28.700 140.690 30.700 ;
        RECT 140.950 28.700 141.120 30.700 ;
        RECT 141.380 28.700 141.550 30.700 ;
        RECT 141.810 28.700 141.980 30.700 ;
        RECT 142.240 28.700 142.410 30.700 ;
        RECT 142.670 28.700 142.840 30.700 ;
        RECT 143.100 28.700 143.270 30.700 ;
        RECT 143.530 28.700 143.700 30.700 ;
        RECT 136.040 28.200 136.570 28.530 ;
        RECT 136.900 28.200 137.430 28.530 ;
        RECT 137.760 28.200 138.290 28.530 ;
        RECT 138.620 28.200 139.150 28.530 ;
        RECT 139.480 28.200 140.010 28.530 ;
        RECT 140.340 28.200 140.870 28.530 ;
        RECT 141.200 28.200 141.730 28.530 ;
        RECT 142.060 28.200 142.590 28.530 ;
        RECT 142.920 28.200 143.450 28.530 ;
        RECT 144.200 27.730 144.370 31.160 ;
        RECT 64.700 23.590 94.610 23.760 ;
        RECT 124.810 22.645 124.980 25.330 ;
        RECT 125.730 24.615 126.260 24.945 ;
        RECT 126.590 24.615 127.120 24.945 ;
        RECT 127.450 24.615 127.980 24.945 ;
        RECT 128.310 24.615 128.840 24.945 ;
        RECT 125.480 23.445 125.650 24.445 ;
        RECT 125.910 23.445 126.080 24.445 ;
        RECT 126.340 23.445 126.510 24.445 ;
        RECT 126.770 23.445 126.940 24.445 ;
        RECT 127.200 23.445 127.370 24.445 ;
        RECT 127.630 23.445 127.800 24.445 ;
        RECT 128.060 23.445 128.230 24.445 ;
        RECT 128.490 23.445 128.660 24.445 ;
        RECT 128.920 23.445 129.090 24.445 ;
        RECT 125.730 22.945 126.260 23.275 ;
        RECT 126.590 22.945 127.120 23.275 ;
        RECT 127.450 22.945 127.980 23.275 ;
        RECT 128.310 22.945 128.840 23.275 ;
        RECT 129.590 22.645 129.760 25.330 ;
        RECT 135.120 24.915 135.290 27.320 ;
        RECT 136.040 26.520 136.570 26.850 ;
        RECT 136.900 26.520 137.430 26.850 ;
        RECT 137.760 26.520 138.290 26.850 ;
        RECT 138.620 26.520 139.150 26.850 ;
        RECT 139.480 26.520 140.010 26.850 ;
        RECT 140.340 26.520 140.870 26.850 ;
        RECT 141.200 26.520 141.730 26.850 ;
        RECT 142.060 26.520 142.590 26.850 ;
        RECT 142.920 26.520 143.450 26.850 ;
        RECT 135.790 25.350 135.960 26.350 ;
        RECT 136.220 25.350 136.390 26.350 ;
        RECT 136.650 25.350 136.820 26.350 ;
        RECT 137.080 25.350 137.250 26.350 ;
        RECT 137.510 25.350 137.680 26.350 ;
        RECT 137.940 25.350 138.110 26.350 ;
        RECT 138.370 25.350 138.540 26.350 ;
        RECT 138.800 25.350 138.970 26.350 ;
        RECT 139.230 25.350 139.400 26.350 ;
        RECT 139.660 25.350 139.830 26.350 ;
        RECT 140.090 25.350 140.260 26.350 ;
        RECT 140.520 25.350 140.690 26.350 ;
        RECT 140.950 25.350 141.120 26.350 ;
        RECT 141.380 25.350 141.550 26.350 ;
        RECT 141.810 25.350 141.980 26.350 ;
        RECT 142.240 25.350 142.410 26.350 ;
        RECT 142.670 25.350 142.840 26.350 ;
        RECT 143.100 25.350 143.270 26.350 ;
        RECT 143.530 25.350 143.700 26.350 ;
        RECT 144.200 24.915 144.370 27.320 ;
        RECT 135.120 24.745 144.370 24.915 ;
        RECT 124.810 22.475 129.760 22.645 ;
        RECT 135.120 22.140 144.370 22.310 ;
        RECT 69.190 21.960 90.060 22.130 ;
        RECT 69.190 19.360 69.360 21.960 ;
        RECT 70.245 21.330 72.215 21.660 ;
        RECT 72.840 21.330 74.450 21.660 ;
        RECT 75.120 21.330 76.730 21.660 ;
        RECT 77.365 21.330 79.335 21.660 ;
        RECT 79.925 21.330 81.895 21.660 ;
        RECT 82.520 21.330 84.130 21.660 ;
        RECT 84.800 21.330 86.410 21.660 ;
        RECT 87.045 21.330 89.015 21.660 ;
        RECT 69.860 20.160 70.030 21.160 ;
        RECT 71.140 20.160 71.310 21.160 ;
        RECT 72.420 20.160 72.590 21.160 ;
        RECT 74.700 20.160 74.870 21.160 ;
        RECT 76.980 20.160 77.150 21.160 ;
        RECT 78.260 20.160 78.430 21.160 ;
        RECT 79.540 20.160 79.710 21.160 ;
        RECT 80.820 20.160 80.990 21.160 ;
        RECT 82.100 20.160 82.270 21.160 ;
        RECT 84.380 20.160 84.550 21.160 ;
        RECT 86.660 20.160 86.830 21.160 ;
        RECT 87.940 20.160 88.110 21.160 ;
        RECT 89.220 20.160 89.390 21.160 ;
        RECT 70.245 19.660 72.215 19.990 ;
        RECT 72.840 19.660 74.450 19.990 ;
        RECT 75.120 19.660 76.730 19.990 ;
        RECT 77.365 19.660 79.335 19.990 ;
        RECT 79.925 19.660 81.895 19.990 ;
        RECT 87.045 19.660 89.015 19.990 ;
        RECT 89.890 19.360 90.060 21.960 ;
        RECT 69.190 19.190 90.060 19.360 ;
        RECT 94.140 21.075 118.450 21.245 ;
        RECT 94.140 18.670 94.310 21.075 ;
        RECT 94.810 20.115 94.980 20.615 ;
        RECT 97.090 20.115 97.260 20.615 ;
        RECT 99.370 20.115 99.540 20.615 ;
        RECT 101.650 20.115 101.820 20.615 ;
        RECT 103.930 20.115 104.100 20.615 ;
        RECT 106.210 20.115 106.380 20.615 ;
        RECT 108.490 20.115 108.660 20.615 ;
        RECT 110.770 20.115 110.940 20.615 ;
        RECT 113.050 20.115 113.220 20.615 ;
        RECT 115.330 20.115 115.500 20.615 ;
        RECT 117.610 20.115 117.780 20.615 ;
        RECT 95.230 19.615 96.840 19.945 ;
        RECT 97.510 19.615 99.120 19.945 ;
        RECT 99.790 19.615 101.400 19.945 ;
        RECT 102.070 19.615 103.680 19.945 ;
        RECT 104.350 19.615 105.960 19.945 ;
        RECT 106.630 19.615 108.240 19.945 ;
        RECT 108.910 19.615 110.520 19.945 ;
        RECT 111.190 19.615 112.800 19.945 ;
        RECT 113.470 19.615 115.080 19.945 ;
        RECT 115.750 19.615 117.360 19.945 ;
        RECT 118.280 18.670 118.450 21.075 ;
        RECT 135.120 18.710 135.290 22.140 ;
        RECT 135.790 19.680 135.960 21.680 ;
        RECT 136.220 19.680 136.390 21.680 ;
        RECT 136.650 19.680 136.820 21.680 ;
        RECT 137.080 19.680 137.250 21.680 ;
        RECT 137.510 19.680 137.680 21.680 ;
        RECT 137.940 19.680 138.110 21.680 ;
        RECT 138.370 19.680 138.540 21.680 ;
        RECT 138.800 19.680 138.970 21.680 ;
        RECT 139.230 19.680 139.400 21.680 ;
        RECT 139.660 19.680 139.830 21.680 ;
        RECT 140.090 19.680 140.260 21.680 ;
        RECT 140.520 19.680 140.690 21.680 ;
        RECT 140.950 19.680 141.120 21.680 ;
        RECT 141.380 19.680 141.550 21.680 ;
        RECT 141.810 19.680 141.980 21.680 ;
        RECT 142.240 19.680 142.410 21.680 ;
        RECT 142.670 19.680 142.840 21.680 ;
        RECT 143.100 19.680 143.270 21.680 ;
        RECT 143.530 19.680 143.700 21.680 ;
        RECT 136.040 19.180 136.570 19.510 ;
        RECT 136.900 19.180 137.430 19.510 ;
        RECT 137.760 19.180 138.290 19.510 ;
        RECT 138.620 19.180 139.150 19.510 ;
        RECT 139.480 19.180 140.010 19.510 ;
        RECT 140.340 19.180 140.870 19.510 ;
        RECT 141.200 19.180 141.730 19.510 ;
        RECT 142.060 19.180 142.590 19.510 ;
        RECT 142.920 19.180 143.450 19.510 ;
        RECT 144.200 18.710 144.370 22.140 ;
        RECT 55.980 17.705 65.170 17.875 ;
        RECT 55.980 15.605 56.150 17.705 ;
        RECT 57.070 17.075 57.960 17.405 ;
        RECT 63.190 17.075 64.080 17.405 ;
        RECT 56.650 16.405 56.820 16.905 ;
        RECT 57.430 16.405 57.600 16.905 ;
        RECT 58.210 16.405 58.380 16.905 ;
        RECT 60.490 16.405 60.660 16.905 ;
        RECT 62.770 16.405 62.940 16.905 ;
        RECT 63.550 16.405 63.720 16.905 ;
        RECT 64.330 16.405 64.500 16.905 ;
        RECT 58.630 15.905 60.240 16.235 ;
        RECT 60.910 15.905 62.520 16.235 ;
        RECT 65.000 15.605 65.170 17.705 ;
        RECT 55.980 15.435 65.170 15.605 ;
        RECT 69.190 17.705 90.060 17.875 ;
        RECT 69.190 15.605 69.360 17.705 ;
        RECT 70.245 17.075 72.215 17.405 ;
        RECT 72.840 17.075 74.450 17.405 ;
        RECT 75.120 17.075 76.730 17.405 ;
        RECT 77.365 17.075 79.335 17.405 ;
        RECT 79.925 17.075 81.895 17.405 ;
        RECT 87.045 17.075 89.015 17.405 ;
        RECT 69.860 16.405 70.030 16.905 ;
        RECT 71.140 16.405 71.310 16.905 ;
        RECT 72.420 16.405 72.590 16.905 ;
        RECT 74.700 16.405 74.870 16.905 ;
        RECT 76.980 16.405 77.150 16.905 ;
        RECT 78.260 16.405 78.430 16.905 ;
        RECT 79.540 16.405 79.710 16.905 ;
        RECT 80.820 16.405 80.990 16.905 ;
        RECT 82.100 16.405 82.270 16.905 ;
        RECT 84.380 16.405 84.550 16.905 ;
        RECT 86.660 16.405 86.830 16.905 ;
        RECT 87.940 16.405 88.110 16.905 ;
        RECT 89.220 16.405 89.390 16.905 ;
        RECT 70.245 15.905 72.215 16.235 ;
        RECT 72.840 15.905 74.450 16.235 ;
        RECT 75.120 15.905 76.730 16.235 ;
        RECT 77.365 15.905 79.335 16.235 ;
        RECT 79.925 15.905 81.895 16.235 ;
        RECT 82.520 15.905 84.130 16.235 ;
        RECT 84.800 15.905 86.410 16.235 ;
        RECT 87.045 15.905 89.015 16.235 ;
        RECT 89.890 15.605 90.060 17.705 ;
        RECT 69.190 15.435 90.060 15.605 ;
        RECT 94.140 14.855 94.310 18.285 ;
        RECT 95.230 16.485 96.840 16.815 ;
        RECT 97.510 16.485 99.120 16.815 ;
        RECT 99.790 16.485 101.400 16.815 ;
        RECT 102.070 16.485 103.680 16.815 ;
        RECT 104.350 16.485 105.960 16.815 ;
        RECT 106.630 16.485 108.240 16.815 ;
        RECT 108.910 16.485 110.520 16.815 ;
        RECT 111.190 16.485 112.800 16.815 ;
        RECT 113.470 16.485 115.080 16.815 ;
        RECT 115.750 16.485 117.360 16.815 ;
        RECT 94.810 15.315 94.980 16.315 ;
        RECT 97.090 15.315 97.260 16.315 ;
        RECT 99.370 15.315 99.540 16.315 ;
        RECT 101.650 15.315 101.820 16.315 ;
        RECT 103.930 15.315 104.100 16.315 ;
        RECT 106.210 15.315 106.380 16.315 ;
        RECT 108.490 15.315 108.660 16.315 ;
        RECT 110.770 15.315 110.940 16.315 ;
        RECT 113.050 15.315 113.220 16.315 ;
        RECT 115.330 15.315 115.500 16.315 ;
        RECT 117.610 15.315 117.780 16.315 ;
        RECT 118.280 14.855 118.450 18.285 ;
        RECT 135.120 15.895 135.290 18.300 ;
        RECT 136.040 17.500 136.570 17.830 ;
        RECT 136.900 17.500 137.430 17.830 ;
        RECT 137.760 17.500 138.290 17.830 ;
        RECT 138.620 17.500 139.150 17.830 ;
        RECT 139.480 17.500 140.010 17.830 ;
        RECT 140.340 17.500 140.870 17.830 ;
        RECT 141.200 17.500 141.730 17.830 ;
        RECT 142.060 17.500 142.590 17.830 ;
        RECT 142.920 17.500 143.450 17.830 ;
        RECT 135.790 16.330 135.960 17.330 ;
        RECT 136.220 16.330 136.390 17.330 ;
        RECT 136.650 16.330 136.820 17.330 ;
        RECT 137.080 16.330 137.250 17.330 ;
        RECT 137.510 16.330 137.680 17.330 ;
        RECT 137.940 16.330 138.110 17.330 ;
        RECT 138.370 16.330 138.540 17.330 ;
        RECT 138.800 16.330 138.970 17.330 ;
        RECT 139.230 16.330 139.400 17.330 ;
        RECT 139.660 16.330 139.830 17.330 ;
        RECT 140.090 16.330 140.260 17.330 ;
        RECT 140.520 16.330 140.690 17.330 ;
        RECT 140.950 16.330 141.120 17.330 ;
        RECT 141.380 16.330 141.550 17.330 ;
        RECT 141.810 16.330 141.980 17.330 ;
        RECT 142.240 16.330 142.410 17.330 ;
        RECT 142.670 16.330 142.840 17.330 ;
        RECT 143.100 16.330 143.270 17.330 ;
        RECT 143.530 16.330 143.700 17.330 ;
        RECT 144.200 15.895 144.370 18.300 ;
        RECT 135.120 15.725 144.370 15.895 ;
        RECT 94.140 14.685 118.450 14.855 ;
        RECT 55.980 13.540 95.650 13.710 ;
        RECT 55.980 7.350 56.150 13.540 ;
        RECT 58.630 12.910 60.240 13.240 ;
        RECT 60.910 12.910 62.520 13.240 ;
        RECT 66.310 12.910 67.920 13.240 ;
        RECT 68.590 12.910 70.200 13.240 ;
        RECT 70.870 12.910 72.480 13.240 ;
        RECT 73.150 12.910 74.760 13.240 ;
        RECT 75.430 12.910 77.040 13.240 ;
        RECT 77.710 12.910 79.320 13.240 ;
        RECT 79.990 12.910 81.600 13.240 ;
        RECT 82.270 12.910 83.880 13.240 ;
        RECT 84.550 12.910 86.160 13.240 ;
        RECT 86.830 12.910 88.440 13.240 ;
        RECT 89.110 12.910 90.720 13.240 ;
        RECT 91.390 12.910 93.000 13.240 ;
        RECT 56.650 11.740 56.820 12.740 ;
        RECT 57.430 11.740 57.600 12.740 ;
        RECT 58.210 11.740 58.380 12.740 ;
        RECT 60.490 11.740 60.660 12.740 ;
        RECT 62.770 11.740 62.940 12.740 ;
        RECT 63.550 11.740 63.720 12.740 ;
        RECT 64.330 11.740 64.500 12.740 ;
        RECT 65.110 11.740 65.280 12.740 ;
        RECT 65.890 11.740 66.060 12.740 ;
        RECT 68.170 11.740 68.340 12.740 ;
        RECT 70.450 11.740 70.620 12.740 ;
        RECT 72.730 11.740 72.900 12.740 ;
        RECT 75.010 11.740 75.180 12.740 ;
        RECT 77.290 11.740 77.460 12.740 ;
        RECT 79.570 11.740 79.740 12.740 ;
        RECT 81.850 11.740 82.020 12.740 ;
        RECT 84.130 11.740 84.300 12.740 ;
        RECT 86.410 11.740 86.580 12.740 ;
        RECT 88.690 11.740 88.860 12.740 ;
        RECT 90.970 11.740 91.140 12.740 ;
        RECT 93.250 11.740 93.420 12.740 ;
        RECT 94.030 11.740 94.200 12.740 ;
        RECT 94.810 11.740 94.980 12.740 ;
        RECT 57.070 11.240 57.960 11.570 ;
        RECT 63.190 11.240 64.080 11.570 ;
        RECT 64.750 11.240 65.640 11.570 ;
        RECT 66.310 11.240 67.920 11.570 ;
        RECT 68.590 11.240 70.200 11.570 ;
        RECT 70.870 11.240 72.480 11.570 ;
        RECT 73.150 11.240 74.760 11.570 ;
        RECT 75.430 11.240 77.040 11.570 ;
        RECT 77.710 11.240 79.320 11.570 ;
        RECT 79.990 11.240 81.600 11.570 ;
        RECT 82.270 11.240 83.880 11.570 ;
        RECT 84.550 11.240 86.160 11.570 ;
        RECT 86.830 11.240 88.440 11.570 ;
        RECT 89.110 11.240 90.720 11.570 ;
        RECT 91.390 11.240 93.000 11.570 ;
        RECT 93.670 11.240 94.560 11.570 ;
        RECT 66.310 9.320 67.920 9.650 ;
        RECT 68.590 9.320 70.200 9.650 ;
        RECT 70.870 9.320 72.480 9.650 ;
        RECT 73.150 9.320 74.760 9.650 ;
        RECT 75.430 9.320 77.040 9.650 ;
        RECT 82.270 9.320 83.880 9.650 ;
        RECT 84.550 9.320 86.160 9.650 ;
        RECT 86.830 9.320 88.440 9.650 ;
        RECT 89.110 9.320 90.720 9.650 ;
        RECT 91.390 9.320 93.000 9.650 ;
        RECT 65.890 8.150 66.060 9.150 ;
        RECT 68.170 8.150 68.340 9.150 ;
        RECT 70.450 8.150 70.620 9.150 ;
        RECT 72.730 8.150 72.900 9.150 ;
        RECT 75.010 8.150 75.180 9.150 ;
        RECT 77.290 8.150 77.460 9.150 ;
        RECT 79.570 8.150 79.740 9.150 ;
        RECT 81.850 8.150 82.020 9.150 ;
        RECT 84.130 8.150 84.300 9.150 ;
        RECT 86.410 8.150 86.580 9.150 ;
        RECT 88.690 8.150 88.860 9.150 ;
        RECT 90.970 8.150 91.140 9.150 ;
        RECT 93.250 8.150 93.420 9.150 ;
        RECT 77.710 7.650 79.320 7.980 ;
        RECT 79.990 7.650 81.600 7.980 ;
        RECT 95.480 7.350 95.650 13.540 ;
        RECT 55.980 7.180 95.650 7.350 ;
      LAYER mcon ;
        RECT 137.170 77.865 137.340 78.035 ;
        RECT 137.610 77.925 137.780 78.095 ;
        RECT 137.970 77.925 138.140 78.095 ;
        RECT 138.330 77.925 138.500 78.095 ;
        RECT 138.690 77.925 138.860 78.095 ;
        RECT 139.050 77.925 139.220 78.095 ;
        RECT 139.410 77.925 139.580 78.095 ;
        RECT 139.770 77.925 139.940 78.095 ;
        RECT 140.130 77.925 140.300 78.095 ;
        RECT 140.490 77.925 140.660 78.095 ;
        RECT 140.850 77.925 141.020 78.095 ;
        RECT 141.210 77.925 141.380 78.095 ;
        RECT 141.570 77.925 141.740 78.095 ;
        RECT 141.930 77.925 142.100 78.095 ;
        RECT 142.290 77.925 142.460 78.095 ;
        RECT 142.650 77.925 142.820 78.095 ;
        RECT 143.010 77.925 143.180 78.095 ;
        RECT 143.370 77.925 143.540 78.095 ;
        RECT 143.730 77.925 143.900 78.095 ;
        RECT 144.090 77.925 144.260 78.095 ;
        RECT 144.450 77.925 144.620 78.095 ;
        RECT 144.810 77.925 144.980 78.095 ;
        RECT 145.170 77.925 145.340 78.095 ;
        RECT 145.530 77.925 145.700 78.095 ;
        RECT 145.890 77.925 146.060 78.095 ;
        RECT 146.250 77.925 146.420 78.095 ;
        RECT 146.610 77.925 146.780 78.095 ;
        RECT 146.970 77.925 147.140 78.095 ;
        RECT 137.170 77.505 137.340 77.675 ;
        RECT 137.170 77.145 137.340 77.315 ;
        RECT 141.670 77.375 141.840 77.545 ;
        RECT 142.530 77.375 142.700 77.545 ;
        RECT 147.030 77.315 147.200 77.485 ;
        RECT 42.770 76.620 42.940 76.790 ;
        RECT 43.130 76.680 43.300 76.850 ;
        RECT 43.490 76.680 43.660 76.850 ;
        RECT 43.850 76.680 44.020 76.850 ;
        RECT 44.210 76.680 44.380 76.850 ;
        RECT 44.570 76.680 44.740 76.850 ;
        RECT 44.930 76.680 45.100 76.850 ;
        RECT 45.290 76.680 45.460 76.850 ;
        RECT 45.650 76.680 45.820 76.850 ;
        RECT 46.010 76.680 46.180 76.850 ;
        RECT 46.370 76.680 46.540 76.850 ;
        RECT 46.730 76.680 46.900 76.850 ;
        RECT 47.090 76.680 47.260 76.850 ;
        RECT 47.450 76.680 47.620 76.850 ;
        RECT 47.810 76.680 47.980 76.850 ;
        RECT 48.170 76.680 48.340 76.850 ;
        RECT 48.530 76.680 48.700 76.850 ;
        RECT 48.890 76.680 49.060 76.850 ;
        RECT 49.250 76.680 49.420 76.850 ;
        RECT 49.610 76.680 49.780 76.850 ;
        RECT 49.970 76.680 50.140 76.850 ;
        RECT 50.330 76.680 50.500 76.850 ;
        RECT 50.690 76.680 50.860 76.850 ;
        RECT 51.050 76.680 51.220 76.850 ;
        RECT 51.410 76.680 51.580 76.850 ;
        RECT 51.770 76.680 51.940 76.850 ;
        RECT 52.130 76.680 52.300 76.850 ;
        RECT 52.490 76.680 52.660 76.850 ;
        RECT 52.850 76.680 53.020 76.850 ;
        RECT 53.210 76.680 53.380 76.850 ;
        RECT 53.570 76.680 53.740 76.850 ;
        RECT 53.930 76.680 54.100 76.850 ;
        RECT 54.290 76.680 54.460 76.850 ;
        RECT 54.650 76.680 54.820 76.850 ;
        RECT 55.010 76.680 55.180 76.850 ;
        RECT 55.370 76.680 55.540 76.850 ;
        RECT 55.730 76.680 55.900 76.850 ;
        RECT 56.090 76.680 56.260 76.850 ;
        RECT 56.450 76.680 56.620 76.850 ;
        RECT 56.810 76.680 56.980 76.850 ;
        RECT 57.170 76.680 57.340 76.850 ;
        RECT 57.530 76.680 57.700 76.850 ;
        RECT 57.890 76.680 58.060 76.850 ;
        RECT 58.250 76.680 58.420 76.850 ;
        RECT 58.610 76.680 58.780 76.850 ;
        RECT 58.970 76.680 59.140 76.850 ;
        RECT 59.330 76.680 59.500 76.850 ;
        RECT 59.690 76.680 59.860 76.850 ;
        RECT 60.050 76.680 60.220 76.850 ;
        RECT 60.410 76.680 60.580 76.850 ;
        RECT 60.770 76.680 60.940 76.850 ;
        RECT 61.130 76.680 61.300 76.850 ;
        RECT 61.490 76.680 61.660 76.850 ;
        RECT 61.850 76.680 62.020 76.850 ;
        RECT 62.210 76.680 62.380 76.850 ;
        RECT 62.570 76.680 62.740 76.850 ;
        RECT 62.930 76.680 63.100 76.850 ;
        RECT 63.290 76.680 63.460 76.850 ;
        RECT 63.650 76.680 63.820 76.850 ;
        RECT 64.010 76.680 64.180 76.850 ;
        RECT 64.370 76.680 64.540 76.850 ;
        RECT 64.730 76.680 64.900 76.850 ;
        RECT 65.090 76.680 65.260 76.850 ;
        RECT 65.450 76.680 65.620 76.850 ;
        RECT 65.810 76.680 65.980 76.850 ;
        RECT 66.170 76.680 66.340 76.850 ;
        RECT 66.530 76.680 66.700 76.850 ;
        RECT 66.890 76.680 67.060 76.850 ;
        RECT 67.250 76.680 67.420 76.850 ;
        RECT 67.610 76.680 67.780 76.850 ;
        RECT 67.970 76.680 68.140 76.850 ;
        RECT 68.330 76.680 68.500 76.850 ;
        RECT 68.690 76.680 68.860 76.850 ;
        RECT 69.050 76.680 69.220 76.850 ;
        RECT 69.410 76.680 69.580 76.850 ;
        RECT 69.770 76.680 69.940 76.850 ;
        RECT 70.130 76.680 70.300 76.850 ;
        RECT 70.490 76.680 70.660 76.850 ;
        RECT 70.850 76.680 71.020 76.850 ;
        RECT 71.210 76.680 71.380 76.850 ;
        RECT 71.570 76.680 71.740 76.850 ;
        RECT 71.930 76.680 72.100 76.850 ;
        RECT 72.290 76.680 72.460 76.850 ;
        RECT 72.650 76.680 72.820 76.850 ;
        RECT 73.010 76.680 73.180 76.850 ;
        RECT 73.370 76.680 73.540 76.850 ;
        RECT 73.730 76.680 73.900 76.850 ;
        RECT 74.090 76.680 74.260 76.850 ;
        RECT 74.450 76.680 74.620 76.850 ;
        RECT 74.810 76.680 74.980 76.850 ;
        RECT 75.170 76.680 75.340 76.850 ;
        RECT 75.530 76.680 75.700 76.850 ;
        RECT 75.890 76.680 76.060 76.850 ;
        RECT 76.250 76.680 76.420 76.850 ;
        RECT 76.610 76.680 76.780 76.850 ;
        RECT 76.970 76.680 77.140 76.850 ;
        RECT 77.330 76.680 77.500 76.850 ;
        RECT 77.690 76.680 77.860 76.850 ;
        RECT 78.050 76.680 78.220 76.850 ;
        RECT 78.410 76.680 78.580 76.850 ;
        RECT 78.770 76.680 78.940 76.850 ;
        RECT 79.130 76.680 79.300 76.850 ;
        RECT 79.490 76.680 79.660 76.850 ;
        RECT 79.850 76.680 80.020 76.850 ;
        RECT 80.210 76.680 80.380 76.850 ;
        RECT 80.570 76.680 80.740 76.850 ;
        RECT 80.930 76.680 81.100 76.850 ;
        RECT 81.290 76.680 81.460 76.850 ;
        RECT 81.650 76.680 81.820 76.850 ;
        RECT 82.010 76.680 82.180 76.850 ;
        RECT 82.370 76.680 82.540 76.850 ;
        RECT 82.730 76.680 82.900 76.850 ;
        RECT 83.090 76.680 83.260 76.850 ;
        RECT 83.450 76.680 83.620 76.850 ;
        RECT 83.810 76.680 83.980 76.850 ;
        RECT 84.170 76.680 84.340 76.850 ;
        RECT 84.530 76.680 84.700 76.850 ;
        RECT 84.890 76.680 85.060 76.850 ;
        RECT 85.250 76.680 85.420 76.850 ;
        RECT 85.610 76.680 85.780 76.850 ;
        RECT 85.970 76.680 86.140 76.850 ;
        RECT 86.330 76.680 86.500 76.850 ;
        RECT 86.690 76.680 86.860 76.850 ;
        RECT 87.050 76.680 87.220 76.850 ;
        RECT 87.410 76.680 87.580 76.850 ;
        RECT 87.770 76.680 87.940 76.850 ;
        RECT 88.130 76.680 88.300 76.850 ;
        RECT 88.490 76.680 88.660 76.850 ;
        RECT 88.850 76.680 89.020 76.850 ;
        RECT 89.210 76.680 89.380 76.850 ;
        RECT 89.570 76.680 89.740 76.850 ;
        RECT 89.930 76.680 90.100 76.850 ;
        RECT 90.290 76.680 90.460 76.850 ;
        RECT 90.650 76.680 90.820 76.850 ;
        RECT 91.010 76.680 91.180 76.850 ;
        RECT 91.370 76.680 91.540 76.850 ;
        RECT 91.730 76.680 91.900 76.850 ;
        RECT 92.090 76.680 92.260 76.850 ;
        RECT 92.450 76.680 92.620 76.850 ;
        RECT 92.810 76.680 92.980 76.850 ;
        RECT 93.170 76.680 93.340 76.850 ;
        RECT 93.530 76.680 93.700 76.850 ;
        RECT 93.890 76.680 94.060 76.850 ;
        RECT 94.250 76.680 94.420 76.850 ;
        RECT 94.610 76.680 94.780 76.850 ;
        RECT 94.970 76.680 95.140 76.850 ;
        RECT 95.330 76.680 95.500 76.850 ;
        RECT 95.690 76.680 95.860 76.850 ;
        RECT 96.050 76.680 96.220 76.850 ;
        RECT 96.410 76.680 96.580 76.850 ;
        RECT 96.770 76.680 96.940 76.850 ;
        RECT 97.130 76.680 97.300 76.850 ;
        RECT 97.490 76.680 97.660 76.850 ;
        RECT 97.850 76.680 98.020 76.850 ;
        RECT 98.210 76.680 98.380 76.850 ;
        RECT 98.570 76.680 98.740 76.850 ;
        RECT 98.930 76.680 99.100 76.850 ;
        RECT 99.290 76.680 99.460 76.850 ;
        RECT 99.650 76.680 99.820 76.850 ;
        RECT 100.010 76.680 100.180 76.850 ;
        RECT 100.370 76.680 100.540 76.850 ;
        RECT 100.730 76.680 100.900 76.850 ;
        RECT 101.090 76.680 101.260 76.850 ;
        RECT 101.450 76.680 101.620 76.850 ;
        RECT 101.810 76.680 101.980 76.850 ;
        RECT 102.170 76.680 102.340 76.850 ;
        RECT 102.530 76.680 102.700 76.850 ;
        RECT 102.890 76.680 103.060 76.850 ;
        RECT 103.250 76.680 103.420 76.850 ;
        RECT 103.610 76.680 103.780 76.850 ;
        RECT 103.970 76.680 104.140 76.850 ;
        RECT 104.330 76.680 104.500 76.850 ;
        RECT 104.690 76.680 104.860 76.850 ;
        RECT 105.050 76.680 105.220 76.850 ;
        RECT 105.410 76.680 105.580 76.850 ;
        RECT 105.770 76.680 105.940 76.850 ;
        RECT 106.130 76.680 106.300 76.850 ;
        RECT 106.490 76.680 106.660 76.850 ;
        RECT 106.850 76.680 107.020 76.850 ;
        RECT 107.210 76.680 107.380 76.850 ;
        RECT 107.570 76.680 107.740 76.850 ;
        RECT 107.930 76.680 108.100 76.850 ;
        RECT 108.290 76.680 108.460 76.850 ;
        RECT 108.650 76.680 108.820 76.850 ;
        RECT 109.010 76.680 109.180 76.850 ;
        RECT 109.370 76.680 109.540 76.850 ;
        RECT 109.730 76.680 109.900 76.850 ;
        RECT 110.090 76.680 110.260 76.850 ;
        RECT 110.450 76.680 110.620 76.850 ;
        RECT 110.810 76.680 110.980 76.850 ;
        RECT 111.170 76.680 111.340 76.850 ;
        RECT 111.530 76.680 111.700 76.850 ;
        RECT 111.890 76.680 112.060 76.850 ;
        RECT 112.250 76.680 112.420 76.850 ;
        RECT 112.610 76.680 112.780 76.850 ;
        RECT 112.970 76.680 113.140 76.850 ;
        RECT 113.330 76.680 113.500 76.850 ;
        RECT 113.690 76.680 113.860 76.850 ;
        RECT 114.050 76.680 114.220 76.850 ;
        RECT 114.410 76.680 114.580 76.850 ;
        RECT 114.770 76.680 114.940 76.850 ;
        RECT 115.130 76.680 115.300 76.850 ;
        RECT 115.490 76.680 115.660 76.850 ;
        RECT 115.850 76.680 116.020 76.850 ;
        RECT 116.210 76.680 116.380 76.850 ;
        RECT 116.570 76.680 116.740 76.850 ;
        RECT 116.930 76.680 117.100 76.850 ;
        RECT 117.290 76.680 117.460 76.850 ;
        RECT 117.650 76.680 117.820 76.850 ;
        RECT 118.010 76.680 118.180 76.850 ;
        RECT 118.370 76.680 118.540 76.850 ;
        RECT 118.730 76.680 118.900 76.850 ;
        RECT 119.090 76.680 119.260 76.850 ;
        RECT 119.450 76.680 119.620 76.850 ;
        RECT 119.810 76.680 119.980 76.850 ;
        RECT 120.170 76.680 120.340 76.850 ;
        RECT 120.530 76.680 120.700 76.850 ;
        RECT 120.890 76.680 121.060 76.850 ;
        RECT 121.250 76.680 121.420 76.850 ;
        RECT 121.610 76.680 121.780 76.850 ;
        RECT 121.970 76.680 122.140 76.850 ;
        RECT 122.330 76.680 122.500 76.850 ;
        RECT 122.690 76.680 122.860 76.850 ;
        RECT 123.050 76.680 123.220 76.850 ;
        RECT 123.410 76.680 123.580 76.850 ;
        RECT 123.770 76.680 123.940 76.850 ;
        RECT 124.130 76.680 124.300 76.850 ;
        RECT 124.490 76.680 124.660 76.850 ;
        RECT 124.850 76.680 125.020 76.850 ;
        RECT 125.210 76.680 125.380 76.850 ;
        RECT 125.570 76.680 125.740 76.850 ;
        RECT 125.930 76.680 126.100 76.850 ;
        RECT 126.290 76.680 126.460 76.850 ;
        RECT 126.650 76.680 126.820 76.850 ;
        RECT 127.010 76.680 127.180 76.850 ;
        RECT 127.370 76.680 127.540 76.850 ;
        RECT 127.730 76.680 127.900 76.850 ;
        RECT 128.090 76.680 128.260 76.850 ;
        RECT 128.450 76.680 128.620 76.850 ;
        RECT 128.810 76.680 128.980 76.850 ;
        RECT 129.170 76.680 129.340 76.850 ;
        RECT 129.530 76.680 129.700 76.850 ;
        RECT 129.890 76.680 130.060 76.850 ;
        RECT 130.250 76.680 130.420 76.850 ;
        RECT 130.610 76.680 130.780 76.850 ;
        RECT 42.770 76.260 42.940 76.430 ;
        RECT 42.770 75.900 42.940 76.070 ;
        RECT 43.820 76.130 43.990 76.300 ;
        RECT 44.180 76.130 44.350 76.300 ;
        RECT 44.540 76.130 44.710 76.300 ;
        RECT 44.900 76.130 45.070 76.300 ;
        RECT 45.260 76.130 45.430 76.300 ;
        RECT 46.100 76.130 46.270 76.300 ;
        RECT 46.460 76.130 46.630 76.300 ;
        RECT 46.820 76.130 46.990 76.300 ;
        RECT 47.180 76.130 47.350 76.300 ;
        RECT 47.540 76.130 47.710 76.300 ;
        RECT 48.380 76.130 48.550 76.300 ;
        RECT 48.740 76.130 48.910 76.300 ;
        RECT 49.100 76.130 49.270 76.300 ;
        RECT 49.460 76.130 49.630 76.300 ;
        RECT 49.820 76.130 49.990 76.300 ;
        RECT 50.660 76.130 50.830 76.300 ;
        RECT 51.020 76.130 51.190 76.300 ;
        RECT 51.380 76.130 51.550 76.300 ;
        RECT 51.740 76.130 51.910 76.300 ;
        RECT 52.100 76.130 52.270 76.300 ;
        RECT 52.940 76.130 53.110 76.300 ;
        RECT 53.300 76.130 53.470 76.300 ;
        RECT 53.660 76.130 53.830 76.300 ;
        RECT 54.020 76.130 54.190 76.300 ;
        RECT 54.380 76.130 54.550 76.300 ;
        RECT 55.220 76.130 55.390 76.300 ;
        RECT 55.580 76.130 55.750 76.300 ;
        RECT 55.940 76.130 56.110 76.300 ;
        RECT 56.300 76.130 56.470 76.300 ;
        RECT 56.660 76.130 56.830 76.300 ;
        RECT 57.500 76.130 57.670 76.300 ;
        RECT 57.860 76.130 58.030 76.300 ;
        RECT 58.220 76.130 58.390 76.300 ;
        RECT 58.580 76.130 58.750 76.300 ;
        RECT 58.940 76.130 59.110 76.300 ;
        RECT 59.780 76.130 59.950 76.300 ;
        RECT 60.140 76.130 60.310 76.300 ;
        RECT 60.500 76.130 60.670 76.300 ;
        RECT 60.860 76.130 61.030 76.300 ;
        RECT 61.220 76.130 61.390 76.300 ;
        RECT 62.060 76.130 62.230 76.300 ;
        RECT 62.420 76.130 62.590 76.300 ;
        RECT 62.780 76.130 62.950 76.300 ;
        RECT 63.140 76.130 63.310 76.300 ;
        RECT 63.500 76.130 63.670 76.300 ;
        RECT 64.340 76.130 64.510 76.300 ;
        RECT 64.700 76.130 64.870 76.300 ;
        RECT 65.060 76.130 65.230 76.300 ;
        RECT 65.420 76.130 65.590 76.300 ;
        RECT 65.780 76.130 65.950 76.300 ;
        RECT 66.620 76.130 66.790 76.300 ;
        RECT 66.980 76.130 67.150 76.300 ;
        RECT 67.340 76.130 67.510 76.300 ;
        RECT 67.700 76.130 67.870 76.300 ;
        RECT 68.060 76.130 68.230 76.300 ;
        RECT 68.900 76.130 69.070 76.300 ;
        RECT 69.260 76.130 69.430 76.300 ;
        RECT 69.620 76.130 69.790 76.300 ;
        RECT 69.980 76.130 70.150 76.300 ;
        RECT 70.340 76.130 70.510 76.300 ;
        RECT 71.180 76.130 71.350 76.300 ;
        RECT 71.540 76.130 71.710 76.300 ;
        RECT 71.900 76.130 72.070 76.300 ;
        RECT 72.260 76.130 72.430 76.300 ;
        RECT 72.620 76.130 72.790 76.300 ;
        RECT 73.460 76.130 73.630 76.300 ;
        RECT 73.820 76.130 73.990 76.300 ;
        RECT 74.180 76.130 74.350 76.300 ;
        RECT 74.540 76.130 74.710 76.300 ;
        RECT 74.900 76.130 75.070 76.300 ;
        RECT 75.740 76.130 75.910 76.300 ;
        RECT 76.100 76.130 76.270 76.300 ;
        RECT 76.460 76.130 76.630 76.300 ;
        RECT 76.820 76.130 76.990 76.300 ;
        RECT 77.180 76.130 77.350 76.300 ;
        RECT 78.020 76.130 78.190 76.300 ;
        RECT 78.380 76.130 78.550 76.300 ;
        RECT 78.740 76.130 78.910 76.300 ;
        RECT 79.100 76.130 79.270 76.300 ;
        RECT 79.460 76.130 79.630 76.300 ;
        RECT 80.300 76.130 80.470 76.300 ;
        RECT 80.660 76.130 80.830 76.300 ;
        RECT 81.020 76.130 81.190 76.300 ;
        RECT 81.380 76.130 81.550 76.300 ;
        RECT 81.740 76.130 81.910 76.300 ;
        RECT 82.580 76.130 82.750 76.300 ;
        RECT 82.940 76.130 83.110 76.300 ;
        RECT 83.300 76.130 83.470 76.300 ;
        RECT 83.660 76.130 83.830 76.300 ;
        RECT 84.020 76.130 84.190 76.300 ;
        RECT 84.860 76.130 85.030 76.300 ;
        RECT 85.220 76.130 85.390 76.300 ;
        RECT 85.580 76.130 85.750 76.300 ;
        RECT 85.940 76.130 86.110 76.300 ;
        RECT 86.300 76.130 86.470 76.300 ;
        RECT 87.140 76.130 87.310 76.300 ;
        RECT 87.500 76.130 87.670 76.300 ;
        RECT 87.860 76.130 88.030 76.300 ;
        RECT 88.220 76.130 88.390 76.300 ;
        RECT 88.580 76.130 88.750 76.300 ;
        RECT 89.420 76.130 89.590 76.300 ;
        RECT 89.780 76.130 89.950 76.300 ;
        RECT 90.140 76.130 90.310 76.300 ;
        RECT 90.500 76.130 90.670 76.300 ;
        RECT 90.860 76.130 91.030 76.300 ;
        RECT 91.700 76.130 91.870 76.300 ;
        RECT 92.060 76.130 92.230 76.300 ;
        RECT 92.420 76.130 92.590 76.300 ;
        RECT 92.780 76.130 92.950 76.300 ;
        RECT 93.140 76.130 93.310 76.300 ;
        RECT 93.980 76.130 94.150 76.300 ;
        RECT 94.340 76.130 94.510 76.300 ;
        RECT 94.700 76.130 94.870 76.300 ;
        RECT 95.060 76.130 95.230 76.300 ;
        RECT 95.420 76.130 95.590 76.300 ;
        RECT 96.260 76.130 96.430 76.300 ;
        RECT 96.620 76.130 96.790 76.300 ;
        RECT 96.980 76.130 97.150 76.300 ;
        RECT 97.340 76.130 97.510 76.300 ;
        RECT 97.700 76.130 97.870 76.300 ;
        RECT 98.540 76.130 98.710 76.300 ;
        RECT 98.900 76.130 99.070 76.300 ;
        RECT 99.260 76.130 99.430 76.300 ;
        RECT 99.620 76.130 99.790 76.300 ;
        RECT 99.980 76.130 100.150 76.300 ;
        RECT 100.820 76.130 100.990 76.300 ;
        RECT 101.180 76.130 101.350 76.300 ;
        RECT 101.540 76.130 101.710 76.300 ;
        RECT 101.900 76.130 102.070 76.300 ;
        RECT 102.260 76.130 102.430 76.300 ;
        RECT 103.100 76.130 103.270 76.300 ;
        RECT 103.460 76.130 103.630 76.300 ;
        RECT 103.820 76.130 103.990 76.300 ;
        RECT 104.180 76.130 104.350 76.300 ;
        RECT 104.540 76.130 104.710 76.300 ;
        RECT 105.380 76.130 105.550 76.300 ;
        RECT 105.740 76.130 105.910 76.300 ;
        RECT 106.100 76.130 106.270 76.300 ;
        RECT 106.460 76.130 106.630 76.300 ;
        RECT 106.820 76.130 106.990 76.300 ;
        RECT 107.660 76.130 107.830 76.300 ;
        RECT 108.020 76.130 108.190 76.300 ;
        RECT 108.380 76.130 108.550 76.300 ;
        RECT 108.740 76.130 108.910 76.300 ;
        RECT 109.100 76.130 109.270 76.300 ;
        RECT 109.940 76.130 110.110 76.300 ;
        RECT 110.300 76.130 110.470 76.300 ;
        RECT 110.660 76.130 110.830 76.300 ;
        RECT 111.020 76.130 111.190 76.300 ;
        RECT 111.380 76.130 111.550 76.300 ;
        RECT 112.220 76.130 112.390 76.300 ;
        RECT 112.580 76.130 112.750 76.300 ;
        RECT 112.940 76.130 113.110 76.300 ;
        RECT 113.300 76.130 113.470 76.300 ;
        RECT 113.660 76.130 113.830 76.300 ;
        RECT 114.500 76.130 114.670 76.300 ;
        RECT 114.860 76.130 115.030 76.300 ;
        RECT 115.220 76.130 115.390 76.300 ;
        RECT 115.580 76.130 115.750 76.300 ;
        RECT 115.940 76.130 116.110 76.300 ;
        RECT 116.780 76.130 116.950 76.300 ;
        RECT 117.140 76.130 117.310 76.300 ;
        RECT 117.500 76.130 117.670 76.300 ;
        RECT 117.860 76.130 118.030 76.300 ;
        RECT 118.220 76.130 118.390 76.300 ;
        RECT 119.060 76.130 119.230 76.300 ;
        RECT 119.420 76.130 119.590 76.300 ;
        RECT 119.780 76.130 119.950 76.300 ;
        RECT 120.140 76.130 120.310 76.300 ;
        RECT 120.500 76.130 120.670 76.300 ;
        RECT 121.340 76.130 121.510 76.300 ;
        RECT 121.700 76.130 121.870 76.300 ;
        RECT 122.060 76.130 122.230 76.300 ;
        RECT 122.420 76.130 122.590 76.300 ;
        RECT 122.780 76.130 122.950 76.300 ;
        RECT 123.620 76.130 123.790 76.300 ;
        RECT 123.980 76.130 124.150 76.300 ;
        RECT 124.340 76.130 124.510 76.300 ;
        RECT 124.700 76.130 124.870 76.300 ;
        RECT 125.060 76.130 125.230 76.300 ;
        RECT 125.900 76.130 126.070 76.300 ;
        RECT 126.260 76.130 126.430 76.300 ;
        RECT 126.620 76.130 126.790 76.300 ;
        RECT 126.980 76.130 127.150 76.300 ;
        RECT 127.340 76.130 127.510 76.300 ;
        RECT 128.180 76.130 128.350 76.300 ;
        RECT 128.540 76.130 128.710 76.300 ;
        RECT 128.900 76.130 129.070 76.300 ;
        RECT 129.260 76.130 129.430 76.300 ;
        RECT 129.620 76.130 129.790 76.300 ;
        RECT 130.670 76.140 130.840 76.310 ;
        RECT 42.770 75.540 42.940 75.710 ;
        RECT 42.770 75.180 42.940 75.350 ;
        RECT 43.400 75.625 43.570 75.795 ;
        RECT 43.400 75.265 43.570 75.435 ;
        RECT 45.680 75.625 45.850 75.795 ;
        RECT 45.680 75.265 45.850 75.435 ;
        RECT 47.960 75.625 48.130 75.795 ;
        RECT 47.960 75.265 48.130 75.435 ;
        RECT 50.240 75.625 50.410 75.795 ;
        RECT 50.240 75.265 50.410 75.435 ;
        RECT 52.520 75.625 52.690 75.795 ;
        RECT 52.520 75.265 52.690 75.435 ;
        RECT 54.800 75.625 54.970 75.795 ;
        RECT 54.800 75.265 54.970 75.435 ;
        RECT 57.080 75.625 57.250 75.795 ;
        RECT 57.080 75.265 57.250 75.435 ;
        RECT 59.360 75.625 59.530 75.795 ;
        RECT 59.360 75.265 59.530 75.435 ;
        RECT 61.640 75.625 61.810 75.795 ;
        RECT 61.640 75.265 61.810 75.435 ;
        RECT 63.920 75.625 64.090 75.795 ;
        RECT 63.920 75.265 64.090 75.435 ;
        RECT 66.200 75.625 66.370 75.795 ;
        RECT 66.200 75.265 66.370 75.435 ;
        RECT 68.480 75.625 68.650 75.795 ;
        RECT 68.480 75.265 68.650 75.435 ;
        RECT 70.760 75.625 70.930 75.795 ;
        RECT 70.760 75.265 70.930 75.435 ;
        RECT 73.040 75.625 73.210 75.795 ;
        RECT 73.040 75.265 73.210 75.435 ;
        RECT 75.320 75.625 75.490 75.795 ;
        RECT 75.320 75.265 75.490 75.435 ;
        RECT 77.600 75.625 77.770 75.795 ;
        RECT 77.600 75.265 77.770 75.435 ;
        RECT 79.880 75.625 80.050 75.795 ;
        RECT 79.880 75.265 80.050 75.435 ;
        RECT 82.160 75.625 82.330 75.795 ;
        RECT 82.160 75.265 82.330 75.435 ;
        RECT 84.440 75.625 84.610 75.795 ;
        RECT 84.440 75.265 84.610 75.435 ;
        RECT 86.720 75.625 86.890 75.795 ;
        RECT 86.720 75.265 86.890 75.435 ;
        RECT 89.000 75.625 89.170 75.795 ;
        RECT 89.000 75.265 89.170 75.435 ;
        RECT 91.280 75.625 91.450 75.795 ;
        RECT 91.280 75.265 91.450 75.435 ;
        RECT 93.560 75.625 93.730 75.795 ;
        RECT 93.560 75.265 93.730 75.435 ;
        RECT 95.840 75.625 96.010 75.795 ;
        RECT 95.840 75.265 96.010 75.435 ;
        RECT 98.120 75.625 98.290 75.795 ;
        RECT 98.120 75.265 98.290 75.435 ;
        RECT 100.400 75.625 100.570 75.795 ;
        RECT 100.400 75.265 100.570 75.435 ;
        RECT 102.680 75.625 102.850 75.795 ;
        RECT 102.680 75.265 102.850 75.435 ;
        RECT 104.960 75.625 105.130 75.795 ;
        RECT 104.960 75.265 105.130 75.435 ;
        RECT 107.240 75.625 107.410 75.795 ;
        RECT 107.240 75.265 107.410 75.435 ;
        RECT 109.520 75.625 109.690 75.795 ;
        RECT 109.520 75.265 109.690 75.435 ;
        RECT 111.800 75.625 111.970 75.795 ;
        RECT 111.800 75.265 111.970 75.435 ;
        RECT 114.080 75.625 114.250 75.795 ;
        RECT 114.080 75.265 114.250 75.435 ;
        RECT 116.360 75.625 116.530 75.795 ;
        RECT 116.360 75.265 116.530 75.435 ;
        RECT 118.640 75.625 118.810 75.795 ;
        RECT 118.640 75.265 118.810 75.435 ;
        RECT 120.920 75.625 121.090 75.795 ;
        RECT 120.920 75.265 121.090 75.435 ;
        RECT 123.200 75.625 123.370 75.795 ;
        RECT 123.200 75.265 123.370 75.435 ;
        RECT 125.480 75.625 125.650 75.795 ;
        RECT 125.480 75.265 125.650 75.435 ;
        RECT 127.760 75.625 127.930 75.795 ;
        RECT 127.760 75.265 127.930 75.435 ;
        RECT 130.040 75.625 130.210 75.795 ;
        RECT 130.040 75.265 130.210 75.435 ;
        RECT 130.670 75.780 130.840 75.950 ;
        RECT 130.670 75.420 130.840 75.590 ;
        RECT 137.170 76.785 137.340 76.955 ;
        RECT 137.170 76.425 137.340 76.595 ;
        RECT 137.800 76.870 137.970 77.040 ;
        RECT 137.800 76.510 137.970 76.680 ;
        RECT 138.230 76.870 138.400 77.040 ;
        RECT 138.230 76.510 138.400 76.680 ;
        RECT 138.660 76.870 138.830 77.040 ;
        RECT 138.660 76.510 138.830 76.680 ;
        RECT 139.090 76.870 139.260 77.040 ;
        RECT 139.090 76.510 139.260 76.680 ;
        RECT 139.520 76.870 139.690 77.040 ;
        RECT 139.520 76.510 139.690 76.680 ;
        RECT 139.950 76.870 140.120 77.040 ;
        RECT 139.950 76.510 140.120 76.680 ;
        RECT 140.380 76.870 140.550 77.040 ;
        RECT 140.380 76.510 140.550 76.680 ;
        RECT 140.810 76.870 140.980 77.040 ;
        RECT 140.810 76.510 140.980 76.680 ;
        RECT 141.240 76.870 141.410 77.040 ;
        RECT 141.240 76.510 141.410 76.680 ;
        RECT 141.670 76.870 141.840 77.040 ;
        RECT 141.670 76.510 141.840 76.680 ;
        RECT 142.100 76.870 142.270 77.040 ;
        RECT 142.100 76.510 142.270 76.680 ;
        RECT 142.530 76.870 142.700 77.040 ;
        RECT 142.530 76.510 142.700 76.680 ;
        RECT 142.960 76.870 143.130 77.040 ;
        RECT 142.960 76.510 143.130 76.680 ;
        RECT 143.390 76.870 143.560 77.040 ;
        RECT 143.390 76.510 143.560 76.680 ;
        RECT 143.820 76.870 143.990 77.040 ;
        RECT 143.820 76.510 143.990 76.680 ;
        RECT 144.250 76.870 144.420 77.040 ;
        RECT 144.250 76.510 144.420 76.680 ;
        RECT 144.680 76.870 144.850 77.040 ;
        RECT 144.680 76.510 144.850 76.680 ;
        RECT 145.110 76.870 145.280 77.040 ;
        RECT 145.110 76.510 145.280 76.680 ;
        RECT 145.540 76.870 145.710 77.040 ;
        RECT 145.540 76.510 145.710 76.680 ;
        RECT 145.970 76.870 146.140 77.040 ;
        RECT 145.970 76.510 146.140 76.680 ;
        RECT 146.400 76.870 146.570 77.040 ;
        RECT 146.400 76.510 146.570 76.680 ;
        RECT 147.030 76.955 147.200 77.125 ;
        RECT 147.030 76.595 147.200 76.765 ;
        RECT 137.170 76.065 137.340 76.235 ;
        RECT 138.230 76.005 138.400 76.175 ;
        RECT 139.090 76.005 139.260 76.175 ;
        RECT 139.950 76.005 140.120 76.175 ;
        RECT 140.810 76.005 140.980 76.175 ;
        RECT 143.390 76.005 143.560 76.175 ;
        RECT 144.250 76.005 144.420 76.175 ;
        RECT 145.110 76.005 145.280 76.175 ;
        RECT 145.970 76.005 146.140 76.175 ;
        RECT 147.030 76.235 147.200 76.405 ;
        RECT 147.030 75.875 147.200 76.045 ;
        RECT 137.230 75.455 137.400 75.625 ;
        RECT 137.590 75.455 137.760 75.625 ;
        RECT 137.950 75.455 138.120 75.625 ;
        RECT 138.310 75.455 138.480 75.625 ;
        RECT 138.670 75.455 138.840 75.625 ;
        RECT 139.030 75.455 139.200 75.625 ;
        RECT 139.390 75.455 139.560 75.625 ;
        RECT 139.750 75.455 139.920 75.625 ;
        RECT 140.110 75.455 140.280 75.625 ;
        RECT 140.470 75.455 140.640 75.625 ;
        RECT 140.830 75.455 141.000 75.625 ;
        RECT 141.190 75.455 141.360 75.625 ;
        RECT 141.550 75.455 141.720 75.625 ;
        RECT 141.910 75.455 142.080 75.625 ;
        RECT 142.280 75.455 142.450 75.625 ;
        RECT 142.640 75.455 142.810 75.625 ;
        RECT 143.000 75.455 143.170 75.625 ;
        RECT 143.360 75.455 143.530 75.625 ;
        RECT 143.720 75.455 143.890 75.625 ;
        RECT 144.080 75.455 144.250 75.625 ;
        RECT 144.440 75.455 144.610 75.625 ;
        RECT 144.800 75.455 144.970 75.625 ;
        RECT 145.160 75.455 145.330 75.625 ;
        RECT 145.520 75.455 145.690 75.625 ;
        RECT 145.880 75.455 146.050 75.625 ;
        RECT 146.240 75.455 146.410 75.625 ;
        RECT 146.600 75.455 146.770 75.625 ;
        RECT 147.030 75.515 147.200 75.685 ;
        RECT 130.670 75.060 130.840 75.230 ;
        RECT 42.770 74.820 42.940 74.990 ;
        RECT 48.380 74.760 48.550 74.930 ;
        RECT 48.740 74.760 48.910 74.930 ;
        RECT 49.100 74.760 49.270 74.930 ;
        RECT 49.460 74.760 49.630 74.930 ;
        RECT 49.820 74.760 49.990 74.930 ;
        RECT 50.660 74.760 50.830 74.930 ;
        RECT 51.020 74.760 51.190 74.930 ;
        RECT 51.380 74.760 51.550 74.930 ;
        RECT 51.740 74.760 51.910 74.930 ;
        RECT 52.100 74.760 52.270 74.930 ;
        RECT 52.940 74.760 53.110 74.930 ;
        RECT 53.300 74.760 53.470 74.930 ;
        RECT 53.660 74.760 53.830 74.930 ;
        RECT 54.020 74.760 54.190 74.930 ;
        RECT 54.380 74.760 54.550 74.930 ;
        RECT 55.220 74.760 55.390 74.930 ;
        RECT 55.580 74.760 55.750 74.930 ;
        RECT 55.940 74.760 56.110 74.930 ;
        RECT 56.300 74.760 56.470 74.930 ;
        RECT 56.660 74.760 56.830 74.930 ;
        RECT 57.500 74.760 57.670 74.930 ;
        RECT 57.860 74.760 58.030 74.930 ;
        RECT 58.220 74.760 58.390 74.930 ;
        RECT 58.580 74.760 58.750 74.930 ;
        RECT 58.940 74.760 59.110 74.930 ;
        RECT 59.780 74.760 59.950 74.930 ;
        RECT 60.140 74.760 60.310 74.930 ;
        RECT 60.500 74.760 60.670 74.930 ;
        RECT 60.860 74.760 61.030 74.930 ;
        RECT 61.220 74.760 61.390 74.930 ;
        RECT 62.060 74.760 62.230 74.930 ;
        RECT 62.420 74.760 62.590 74.930 ;
        RECT 62.780 74.760 62.950 74.930 ;
        RECT 63.140 74.760 63.310 74.930 ;
        RECT 63.500 74.760 63.670 74.930 ;
        RECT 64.340 74.760 64.510 74.930 ;
        RECT 64.700 74.760 64.870 74.930 ;
        RECT 65.060 74.760 65.230 74.930 ;
        RECT 65.420 74.760 65.590 74.930 ;
        RECT 65.780 74.760 65.950 74.930 ;
        RECT 66.620 74.760 66.790 74.930 ;
        RECT 66.980 74.760 67.150 74.930 ;
        RECT 67.340 74.760 67.510 74.930 ;
        RECT 67.700 74.760 67.870 74.930 ;
        RECT 68.060 74.760 68.230 74.930 ;
        RECT 68.900 74.760 69.070 74.930 ;
        RECT 69.260 74.760 69.430 74.930 ;
        RECT 69.620 74.760 69.790 74.930 ;
        RECT 69.980 74.760 70.150 74.930 ;
        RECT 70.340 74.760 70.510 74.930 ;
        RECT 71.180 74.760 71.350 74.930 ;
        RECT 71.540 74.760 71.710 74.930 ;
        RECT 71.900 74.760 72.070 74.930 ;
        RECT 72.260 74.760 72.430 74.930 ;
        RECT 72.620 74.760 72.790 74.930 ;
        RECT 73.460 74.760 73.630 74.930 ;
        RECT 73.820 74.760 73.990 74.930 ;
        RECT 74.180 74.760 74.350 74.930 ;
        RECT 74.540 74.760 74.710 74.930 ;
        RECT 74.900 74.760 75.070 74.930 ;
        RECT 75.740 74.760 75.910 74.930 ;
        RECT 76.100 74.760 76.270 74.930 ;
        RECT 76.460 74.760 76.630 74.930 ;
        RECT 76.820 74.760 76.990 74.930 ;
        RECT 77.180 74.760 77.350 74.930 ;
        RECT 78.020 74.760 78.190 74.930 ;
        RECT 78.380 74.760 78.550 74.930 ;
        RECT 78.740 74.760 78.910 74.930 ;
        RECT 79.100 74.760 79.270 74.930 ;
        RECT 79.460 74.760 79.630 74.930 ;
        RECT 80.300 74.760 80.470 74.930 ;
        RECT 80.660 74.760 80.830 74.930 ;
        RECT 81.020 74.760 81.190 74.930 ;
        RECT 81.380 74.760 81.550 74.930 ;
        RECT 81.740 74.760 81.910 74.930 ;
        RECT 82.580 74.760 82.750 74.930 ;
        RECT 82.940 74.760 83.110 74.930 ;
        RECT 83.300 74.760 83.470 74.930 ;
        RECT 83.660 74.760 83.830 74.930 ;
        RECT 84.020 74.760 84.190 74.930 ;
        RECT 84.860 74.760 85.030 74.930 ;
        RECT 85.220 74.760 85.390 74.930 ;
        RECT 85.580 74.760 85.750 74.930 ;
        RECT 85.940 74.760 86.110 74.930 ;
        RECT 86.300 74.760 86.470 74.930 ;
        RECT 87.140 74.760 87.310 74.930 ;
        RECT 87.500 74.760 87.670 74.930 ;
        RECT 87.860 74.760 88.030 74.930 ;
        RECT 88.220 74.760 88.390 74.930 ;
        RECT 88.580 74.760 88.750 74.930 ;
        RECT 89.420 74.760 89.590 74.930 ;
        RECT 89.780 74.760 89.950 74.930 ;
        RECT 90.140 74.760 90.310 74.930 ;
        RECT 90.500 74.760 90.670 74.930 ;
        RECT 90.860 74.760 91.030 74.930 ;
        RECT 91.700 74.760 91.870 74.930 ;
        RECT 92.060 74.760 92.230 74.930 ;
        RECT 92.420 74.760 92.590 74.930 ;
        RECT 92.780 74.760 92.950 74.930 ;
        RECT 93.140 74.760 93.310 74.930 ;
        RECT 93.980 74.760 94.150 74.930 ;
        RECT 94.340 74.760 94.510 74.930 ;
        RECT 94.700 74.760 94.870 74.930 ;
        RECT 95.060 74.760 95.230 74.930 ;
        RECT 95.420 74.760 95.590 74.930 ;
        RECT 96.260 74.760 96.430 74.930 ;
        RECT 96.620 74.760 96.790 74.930 ;
        RECT 96.980 74.760 97.150 74.930 ;
        RECT 97.340 74.760 97.510 74.930 ;
        RECT 97.700 74.760 97.870 74.930 ;
        RECT 98.540 74.760 98.710 74.930 ;
        RECT 98.900 74.760 99.070 74.930 ;
        RECT 99.260 74.760 99.430 74.930 ;
        RECT 99.620 74.760 99.790 74.930 ;
        RECT 99.980 74.760 100.150 74.930 ;
        RECT 100.820 74.760 100.990 74.930 ;
        RECT 101.180 74.760 101.350 74.930 ;
        RECT 101.540 74.760 101.710 74.930 ;
        RECT 101.900 74.760 102.070 74.930 ;
        RECT 102.260 74.760 102.430 74.930 ;
        RECT 103.100 74.760 103.270 74.930 ;
        RECT 103.460 74.760 103.630 74.930 ;
        RECT 103.820 74.760 103.990 74.930 ;
        RECT 104.180 74.760 104.350 74.930 ;
        RECT 104.540 74.760 104.710 74.930 ;
        RECT 105.380 74.760 105.550 74.930 ;
        RECT 105.740 74.760 105.910 74.930 ;
        RECT 106.100 74.760 106.270 74.930 ;
        RECT 106.460 74.760 106.630 74.930 ;
        RECT 106.820 74.760 106.990 74.930 ;
        RECT 107.660 74.760 107.830 74.930 ;
        RECT 108.020 74.760 108.190 74.930 ;
        RECT 108.380 74.760 108.550 74.930 ;
        RECT 108.740 74.760 108.910 74.930 ;
        RECT 109.100 74.760 109.270 74.930 ;
        RECT 109.940 74.760 110.110 74.930 ;
        RECT 110.300 74.760 110.470 74.930 ;
        RECT 110.660 74.760 110.830 74.930 ;
        RECT 111.020 74.760 111.190 74.930 ;
        RECT 111.380 74.760 111.550 74.930 ;
        RECT 112.220 74.760 112.390 74.930 ;
        RECT 112.580 74.760 112.750 74.930 ;
        RECT 112.940 74.760 113.110 74.930 ;
        RECT 113.300 74.760 113.470 74.930 ;
        RECT 113.660 74.760 113.830 74.930 ;
        RECT 114.500 74.760 114.670 74.930 ;
        RECT 114.860 74.760 115.030 74.930 ;
        RECT 115.220 74.760 115.390 74.930 ;
        RECT 115.580 74.760 115.750 74.930 ;
        RECT 115.940 74.760 116.110 74.930 ;
        RECT 128.180 74.760 128.350 74.930 ;
        RECT 128.540 74.760 128.710 74.930 ;
        RECT 128.900 74.760 129.070 74.930 ;
        RECT 129.260 74.760 129.430 74.930 ;
        RECT 129.620 74.760 129.790 74.930 ;
        RECT 130.670 74.700 130.840 74.870 ;
        RECT 42.770 74.460 42.940 74.630 ;
        RECT 42.770 74.100 42.940 74.270 ;
        RECT 42.770 73.740 42.940 73.910 ;
        RECT 43.400 74.255 43.570 74.425 ;
        RECT 43.400 73.895 43.570 74.065 ;
        RECT 45.680 74.255 45.850 74.425 ;
        RECT 45.680 73.895 45.850 74.065 ;
        RECT 47.960 74.255 48.130 74.425 ;
        RECT 47.960 73.895 48.130 74.065 ;
        RECT 50.240 74.255 50.410 74.425 ;
        RECT 50.240 73.895 50.410 74.065 ;
        RECT 52.520 74.255 52.690 74.425 ;
        RECT 52.520 73.895 52.690 74.065 ;
        RECT 54.800 74.255 54.970 74.425 ;
        RECT 54.800 73.895 54.970 74.065 ;
        RECT 57.080 74.255 57.250 74.425 ;
        RECT 57.080 73.895 57.250 74.065 ;
        RECT 59.360 74.255 59.530 74.425 ;
        RECT 59.360 73.895 59.530 74.065 ;
        RECT 61.640 74.255 61.810 74.425 ;
        RECT 61.640 73.895 61.810 74.065 ;
        RECT 63.920 74.255 64.090 74.425 ;
        RECT 63.920 73.895 64.090 74.065 ;
        RECT 66.200 74.255 66.370 74.425 ;
        RECT 66.200 73.895 66.370 74.065 ;
        RECT 68.480 74.255 68.650 74.425 ;
        RECT 68.480 73.895 68.650 74.065 ;
        RECT 70.760 74.255 70.930 74.425 ;
        RECT 70.760 73.895 70.930 74.065 ;
        RECT 73.040 74.255 73.210 74.425 ;
        RECT 73.040 73.895 73.210 74.065 ;
        RECT 75.320 74.255 75.490 74.425 ;
        RECT 75.320 73.895 75.490 74.065 ;
        RECT 77.600 74.255 77.770 74.425 ;
        RECT 77.600 73.895 77.770 74.065 ;
        RECT 79.880 74.255 80.050 74.425 ;
        RECT 79.880 73.895 80.050 74.065 ;
        RECT 82.160 74.255 82.330 74.425 ;
        RECT 82.160 73.895 82.330 74.065 ;
        RECT 84.440 74.255 84.610 74.425 ;
        RECT 84.440 73.895 84.610 74.065 ;
        RECT 86.720 74.255 86.890 74.425 ;
        RECT 86.720 73.895 86.890 74.065 ;
        RECT 89.000 74.255 89.170 74.425 ;
        RECT 89.000 73.895 89.170 74.065 ;
        RECT 91.280 74.255 91.450 74.425 ;
        RECT 91.280 73.895 91.450 74.065 ;
        RECT 93.560 74.255 93.730 74.425 ;
        RECT 93.560 73.895 93.730 74.065 ;
        RECT 95.840 74.255 96.010 74.425 ;
        RECT 95.840 73.895 96.010 74.065 ;
        RECT 98.120 74.255 98.290 74.425 ;
        RECT 98.120 73.895 98.290 74.065 ;
        RECT 100.400 74.255 100.570 74.425 ;
        RECT 100.400 73.895 100.570 74.065 ;
        RECT 102.680 74.255 102.850 74.425 ;
        RECT 102.680 73.895 102.850 74.065 ;
        RECT 104.960 74.255 105.130 74.425 ;
        RECT 104.960 73.895 105.130 74.065 ;
        RECT 107.240 74.255 107.410 74.425 ;
        RECT 107.240 73.895 107.410 74.065 ;
        RECT 109.520 74.255 109.690 74.425 ;
        RECT 109.520 73.895 109.690 74.065 ;
        RECT 111.800 74.255 111.970 74.425 ;
        RECT 111.800 73.895 111.970 74.065 ;
        RECT 114.080 74.255 114.250 74.425 ;
        RECT 114.080 73.895 114.250 74.065 ;
        RECT 116.360 74.255 116.530 74.425 ;
        RECT 116.360 73.895 116.530 74.065 ;
        RECT 118.640 74.255 118.810 74.425 ;
        RECT 118.640 73.895 118.810 74.065 ;
        RECT 120.920 74.255 121.090 74.425 ;
        RECT 120.920 73.895 121.090 74.065 ;
        RECT 123.200 74.255 123.370 74.425 ;
        RECT 123.200 73.895 123.370 74.065 ;
        RECT 125.480 74.255 125.650 74.425 ;
        RECT 125.480 73.895 125.650 74.065 ;
        RECT 127.760 74.255 127.930 74.425 ;
        RECT 127.760 73.895 127.930 74.065 ;
        RECT 130.040 74.255 130.210 74.425 ;
        RECT 130.040 73.895 130.210 74.065 ;
        RECT 130.670 74.340 130.840 74.510 ;
        RECT 130.670 73.980 130.840 74.150 ;
        RECT 42.770 73.380 42.940 73.550 ;
        RECT 43.820 73.390 43.990 73.560 ;
        RECT 44.180 73.390 44.350 73.560 ;
        RECT 44.540 73.390 44.710 73.560 ;
        RECT 44.900 73.390 45.070 73.560 ;
        RECT 45.260 73.390 45.430 73.560 ;
        RECT 46.100 73.390 46.270 73.560 ;
        RECT 46.460 73.390 46.630 73.560 ;
        RECT 46.820 73.390 46.990 73.560 ;
        RECT 47.180 73.390 47.350 73.560 ;
        RECT 47.540 73.390 47.710 73.560 ;
        RECT 48.380 73.390 48.550 73.560 ;
        RECT 48.740 73.390 48.910 73.560 ;
        RECT 49.100 73.390 49.270 73.560 ;
        RECT 49.460 73.390 49.630 73.560 ;
        RECT 49.820 73.390 49.990 73.560 ;
        RECT 50.660 73.390 50.830 73.560 ;
        RECT 51.020 73.390 51.190 73.560 ;
        RECT 51.380 73.390 51.550 73.560 ;
        RECT 51.740 73.390 51.910 73.560 ;
        RECT 52.100 73.390 52.270 73.560 ;
        RECT 52.940 73.390 53.110 73.560 ;
        RECT 53.300 73.390 53.470 73.560 ;
        RECT 53.660 73.390 53.830 73.560 ;
        RECT 54.020 73.390 54.190 73.560 ;
        RECT 54.380 73.390 54.550 73.560 ;
        RECT 55.220 73.390 55.390 73.560 ;
        RECT 55.580 73.390 55.750 73.560 ;
        RECT 55.940 73.390 56.110 73.560 ;
        RECT 56.300 73.390 56.470 73.560 ;
        RECT 56.660 73.390 56.830 73.560 ;
        RECT 57.500 73.390 57.670 73.560 ;
        RECT 57.860 73.390 58.030 73.560 ;
        RECT 58.220 73.390 58.390 73.560 ;
        RECT 58.580 73.390 58.750 73.560 ;
        RECT 58.940 73.390 59.110 73.560 ;
        RECT 59.780 73.390 59.950 73.560 ;
        RECT 60.140 73.390 60.310 73.560 ;
        RECT 60.500 73.390 60.670 73.560 ;
        RECT 60.860 73.390 61.030 73.560 ;
        RECT 61.220 73.390 61.390 73.560 ;
        RECT 62.060 73.390 62.230 73.560 ;
        RECT 62.420 73.390 62.590 73.560 ;
        RECT 62.780 73.390 62.950 73.560 ;
        RECT 63.140 73.390 63.310 73.560 ;
        RECT 63.500 73.390 63.670 73.560 ;
        RECT 64.340 73.390 64.510 73.560 ;
        RECT 64.700 73.390 64.870 73.560 ;
        RECT 65.060 73.390 65.230 73.560 ;
        RECT 65.420 73.390 65.590 73.560 ;
        RECT 65.780 73.390 65.950 73.560 ;
        RECT 66.620 73.390 66.790 73.560 ;
        RECT 66.980 73.390 67.150 73.560 ;
        RECT 67.340 73.390 67.510 73.560 ;
        RECT 67.700 73.390 67.870 73.560 ;
        RECT 68.060 73.390 68.230 73.560 ;
        RECT 68.900 73.390 69.070 73.560 ;
        RECT 69.260 73.390 69.430 73.560 ;
        RECT 69.620 73.390 69.790 73.560 ;
        RECT 69.980 73.390 70.150 73.560 ;
        RECT 70.340 73.390 70.510 73.560 ;
        RECT 71.180 73.390 71.350 73.560 ;
        RECT 71.540 73.390 71.710 73.560 ;
        RECT 71.900 73.390 72.070 73.560 ;
        RECT 72.260 73.390 72.430 73.560 ;
        RECT 72.620 73.390 72.790 73.560 ;
        RECT 73.460 73.390 73.630 73.560 ;
        RECT 73.820 73.390 73.990 73.560 ;
        RECT 74.180 73.390 74.350 73.560 ;
        RECT 74.540 73.390 74.710 73.560 ;
        RECT 74.900 73.390 75.070 73.560 ;
        RECT 75.740 73.390 75.910 73.560 ;
        RECT 76.100 73.390 76.270 73.560 ;
        RECT 76.460 73.390 76.630 73.560 ;
        RECT 76.820 73.390 76.990 73.560 ;
        RECT 77.180 73.390 77.350 73.560 ;
        RECT 78.020 73.390 78.190 73.560 ;
        RECT 78.380 73.390 78.550 73.560 ;
        RECT 78.740 73.390 78.910 73.560 ;
        RECT 79.100 73.390 79.270 73.560 ;
        RECT 79.460 73.390 79.630 73.560 ;
        RECT 80.300 73.390 80.470 73.560 ;
        RECT 80.660 73.390 80.830 73.560 ;
        RECT 81.020 73.390 81.190 73.560 ;
        RECT 81.380 73.390 81.550 73.560 ;
        RECT 81.740 73.390 81.910 73.560 ;
        RECT 82.580 73.390 82.750 73.560 ;
        RECT 82.940 73.390 83.110 73.560 ;
        RECT 83.300 73.390 83.470 73.560 ;
        RECT 83.660 73.390 83.830 73.560 ;
        RECT 84.020 73.390 84.190 73.560 ;
        RECT 84.860 73.390 85.030 73.560 ;
        RECT 85.220 73.390 85.390 73.560 ;
        RECT 85.580 73.390 85.750 73.560 ;
        RECT 85.940 73.390 86.110 73.560 ;
        RECT 86.300 73.390 86.470 73.560 ;
        RECT 87.140 73.390 87.310 73.560 ;
        RECT 87.500 73.390 87.670 73.560 ;
        RECT 87.860 73.390 88.030 73.560 ;
        RECT 88.220 73.390 88.390 73.560 ;
        RECT 88.580 73.390 88.750 73.560 ;
        RECT 89.420 73.390 89.590 73.560 ;
        RECT 89.780 73.390 89.950 73.560 ;
        RECT 90.140 73.390 90.310 73.560 ;
        RECT 90.500 73.390 90.670 73.560 ;
        RECT 90.860 73.390 91.030 73.560 ;
        RECT 91.700 73.390 91.870 73.560 ;
        RECT 92.060 73.390 92.230 73.560 ;
        RECT 92.420 73.390 92.590 73.560 ;
        RECT 92.780 73.390 92.950 73.560 ;
        RECT 93.140 73.390 93.310 73.560 ;
        RECT 93.980 73.390 94.150 73.560 ;
        RECT 94.340 73.390 94.510 73.560 ;
        RECT 94.700 73.390 94.870 73.560 ;
        RECT 95.060 73.390 95.230 73.560 ;
        RECT 95.420 73.390 95.590 73.560 ;
        RECT 96.260 73.390 96.430 73.560 ;
        RECT 96.620 73.390 96.790 73.560 ;
        RECT 96.980 73.390 97.150 73.560 ;
        RECT 97.340 73.390 97.510 73.560 ;
        RECT 97.700 73.390 97.870 73.560 ;
        RECT 98.540 73.390 98.710 73.560 ;
        RECT 98.900 73.390 99.070 73.560 ;
        RECT 99.260 73.390 99.430 73.560 ;
        RECT 99.620 73.390 99.790 73.560 ;
        RECT 99.980 73.390 100.150 73.560 ;
        RECT 100.820 73.390 100.990 73.560 ;
        RECT 101.180 73.390 101.350 73.560 ;
        RECT 101.540 73.390 101.710 73.560 ;
        RECT 101.900 73.390 102.070 73.560 ;
        RECT 102.260 73.390 102.430 73.560 ;
        RECT 103.100 73.390 103.270 73.560 ;
        RECT 103.460 73.390 103.630 73.560 ;
        RECT 103.820 73.390 103.990 73.560 ;
        RECT 104.180 73.390 104.350 73.560 ;
        RECT 104.540 73.390 104.710 73.560 ;
        RECT 105.380 73.390 105.550 73.560 ;
        RECT 105.740 73.390 105.910 73.560 ;
        RECT 106.100 73.390 106.270 73.560 ;
        RECT 106.460 73.390 106.630 73.560 ;
        RECT 106.820 73.390 106.990 73.560 ;
        RECT 107.660 73.390 107.830 73.560 ;
        RECT 108.020 73.390 108.190 73.560 ;
        RECT 108.380 73.390 108.550 73.560 ;
        RECT 108.740 73.390 108.910 73.560 ;
        RECT 109.100 73.390 109.270 73.560 ;
        RECT 109.940 73.390 110.110 73.560 ;
        RECT 110.300 73.390 110.470 73.560 ;
        RECT 110.660 73.390 110.830 73.560 ;
        RECT 111.020 73.390 111.190 73.560 ;
        RECT 111.380 73.390 111.550 73.560 ;
        RECT 112.220 73.390 112.390 73.560 ;
        RECT 112.580 73.390 112.750 73.560 ;
        RECT 112.940 73.390 113.110 73.560 ;
        RECT 113.300 73.390 113.470 73.560 ;
        RECT 113.660 73.390 113.830 73.560 ;
        RECT 114.500 73.390 114.670 73.560 ;
        RECT 114.860 73.390 115.030 73.560 ;
        RECT 115.220 73.390 115.390 73.560 ;
        RECT 115.580 73.390 115.750 73.560 ;
        RECT 115.940 73.390 116.110 73.560 ;
        RECT 116.780 73.390 116.950 73.560 ;
        RECT 117.140 73.390 117.310 73.560 ;
        RECT 117.500 73.390 117.670 73.560 ;
        RECT 117.860 73.390 118.030 73.560 ;
        RECT 118.220 73.390 118.390 73.560 ;
        RECT 119.060 73.390 119.230 73.560 ;
        RECT 119.420 73.390 119.590 73.560 ;
        RECT 119.780 73.390 119.950 73.560 ;
        RECT 120.140 73.390 120.310 73.560 ;
        RECT 120.500 73.390 120.670 73.560 ;
        RECT 121.340 73.390 121.510 73.560 ;
        RECT 121.700 73.390 121.870 73.560 ;
        RECT 122.060 73.390 122.230 73.560 ;
        RECT 122.420 73.390 122.590 73.560 ;
        RECT 122.780 73.390 122.950 73.560 ;
        RECT 123.620 73.390 123.790 73.560 ;
        RECT 123.980 73.390 124.150 73.560 ;
        RECT 124.340 73.390 124.510 73.560 ;
        RECT 124.700 73.390 124.870 73.560 ;
        RECT 125.060 73.390 125.230 73.560 ;
        RECT 125.900 73.390 126.070 73.560 ;
        RECT 126.260 73.390 126.430 73.560 ;
        RECT 126.620 73.390 126.790 73.560 ;
        RECT 126.980 73.390 127.150 73.560 ;
        RECT 127.340 73.390 127.510 73.560 ;
        RECT 128.180 73.390 128.350 73.560 ;
        RECT 128.540 73.390 128.710 73.560 ;
        RECT 128.900 73.390 129.070 73.560 ;
        RECT 129.260 73.390 129.430 73.560 ;
        RECT 129.620 73.390 129.790 73.560 ;
        RECT 130.670 73.620 130.840 73.790 ;
        RECT 130.670 73.260 130.840 73.430 ;
        RECT 42.830 72.840 43.000 73.010 ;
        RECT 43.190 72.840 43.360 73.010 ;
        RECT 43.550 72.840 43.720 73.010 ;
        RECT 43.910 72.840 44.080 73.010 ;
        RECT 44.270 72.840 44.440 73.010 ;
        RECT 44.630 72.840 44.800 73.010 ;
        RECT 44.990 72.840 45.160 73.010 ;
        RECT 45.350 72.840 45.520 73.010 ;
        RECT 45.710 72.840 45.880 73.010 ;
        RECT 46.070 72.840 46.240 73.010 ;
        RECT 46.430 72.840 46.600 73.010 ;
        RECT 46.790 72.840 46.960 73.010 ;
        RECT 47.150 72.840 47.320 73.010 ;
        RECT 47.510 72.840 47.680 73.010 ;
        RECT 47.870 72.840 48.040 73.010 ;
        RECT 48.230 72.840 48.400 73.010 ;
        RECT 48.590 72.840 48.760 73.010 ;
        RECT 48.950 72.840 49.120 73.010 ;
        RECT 49.310 72.840 49.480 73.010 ;
        RECT 49.670 72.840 49.840 73.010 ;
        RECT 50.030 72.840 50.200 73.010 ;
        RECT 50.390 72.840 50.560 73.010 ;
        RECT 50.750 72.840 50.920 73.010 ;
        RECT 51.110 72.840 51.280 73.010 ;
        RECT 51.470 72.840 51.640 73.010 ;
        RECT 51.830 72.840 52.000 73.010 ;
        RECT 52.190 72.840 52.360 73.010 ;
        RECT 52.550 72.840 52.720 73.010 ;
        RECT 52.910 72.840 53.080 73.010 ;
        RECT 53.270 72.840 53.440 73.010 ;
        RECT 53.630 72.840 53.800 73.010 ;
        RECT 53.990 72.840 54.160 73.010 ;
        RECT 54.350 72.840 54.520 73.010 ;
        RECT 54.710 72.840 54.880 73.010 ;
        RECT 55.070 72.840 55.240 73.010 ;
        RECT 55.430 72.840 55.600 73.010 ;
        RECT 55.790 72.840 55.960 73.010 ;
        RECT 56.150 72.840 56.320 73.010 ;
        RECT 56.510 72.840 56.680 73.010 ;
        RECT 56.870 72.840 57.040 73.010 ;
        RECT 57.230 72.840 57.400 73.010 ;
        RECT 57.590 72.840 57.760 73.010 ;
        RECT 57.950 72.840 58.120 73.010 ;
        RECT 58.310 72.840 58.480 73.010 ;
        RECT 58.670 72.840 58.840 73.010 ;
        RECT 59.030 72.840 59.200 73.010 ;
        RECT 59.390 72.840 59.560 73.010 ;
        RECT 59.750 72.840 59.920 73.010 ;
        RECT 60.110 72.840 60.280 73.010 ;
        RECT 60.470 72.840 60.640 73.010 ;
        RECT 60.830 72.840 61.000 73.010 ;
        RECT 61.190 72.840 61.360 73.010 ;
        RECT 61.550 72.840 61.720 73.010 ;
        RECT 61.910 72.840 62.080 73.010 ;
        RECT 62.270 72.840 62.440 73.010 ;
        RECT 62.630 72.840 62.800 73.010 ;
        RECT 62.990 72.840 63.160 73.010 ;
        RECT 63.350 72.840 63.520 73.010 ;
        RECT 63.710 72.840 63.880 73.010 ;
        RECT 64.070 72.840 64.240 73.010 ;
        RECT 64.430 72.840 64.600 73.010 ;
        RECT 64.790 72.840 64.960 73.010 ;
        RECT 65.150 72.840 65.320 73.010 ;
        RECT 65.510 72.840 65.680 73.010 ;
        RECT 65.870 72.840 66.040 73.010 ;
        RECT 66.230 72.840 66.400 73.010 ;
        RECT 66.590 72.840 66.760 73.010 ;
        RECT 66.950 72.840 67.120 73.010 ;
        RECT 67.310 72.840 67.480 73.010 ;
        RECT 67.670 72.840 67.840 73.010 ;
        RECT 68.030 72.840 68.200 73.010 ;
        RECT 68.390 72.840 68.560 73.010 ;
        RECT 68.750 72.840 68.920 73.010 ;
        RECT 69.110 72.840 69.280 73.010 ;
        RECT 69.470 72.840 69.640 73.010 ;
        RECT 69.830 72.840 70.000 73.010 ;
        RECT 70.190 72.840 70.360 73.010 ;
        RECT 70.550 72.840 70.720 73.010 ;
        RECT 70.910 72.840 71.080 73.010 ;
        RECT 71.270 72.840 71.440 73.010 ;
        RECT 71.630 72.840 71.800 73.010 ;
        RECT 71.990 72.840 72.160 73.010 ;
        RECT 72.350 72.840 72.520 73.010 ;
        RECT 72.710 72.840 72.880 73.010 ;
        RECT 73.070 72.840 73.240 73.010 ;
        RECT 73.430 72.840 73.600 73.010 ;
        RECT 73.790 72.840 73.960 73.010 ;
        RECT 74.150 72.840 74.320 73.010 ;
        RECT 74.510 72.840 74.680 73.010 ;
        RECT 74.870 72.840 75.040 73.010 ;
        RECT 75.230 72.840 75.400 73.010 ;
        RECT 75.590 72.840 75.760 73.010 ;
        RECT 75.950 72.840 76.120 73.010 ;
        RECT 76.310 72.840 76.480 73.010 ;
        RECT 76.670 72.840 76.840 73.010 ;
        RECT 77.030 72.840 77.200 73.010 ;
        RECT 77.390 72.840 77.560 73.010 ;
        RECT 77.750 72.840 77.920 73.010 ;
        RECT 78.110 72.840 78.280 73.010 ;
        RECT 78.470 72.840 78.640 73.010 ;
        RECT 78.830 72.840 79.000 73.010 ;
        RECT 79.190 72.840 79.360 73.010 ;
        RECT 79.550 72.840 79.720 73.010 ;
        RECT 79.910 72.840 80.080 73.010 ;
        RECT 80.270 72.840 80.440 73.010 ;
        RECT 80.630 72.840 80.800 73.010 ;
        RECT 80.990 72.840 81.160 73.010 ;
        RECT 81.350 72.840 81.520 73.010 ;
        RECT 81.710 72.840 81.880 73.010 ;
        RECT 82.070 72.840 82.240 73.010 ;
        RECT 82.430 72.840 82.600 73.010 ;
        RECT 82.790 72.840 82.960 73.010 ;
        RECT 83.150 72.840 83.320 73.010 ;
        RECT 83.510 72.840 83.680 73.010 ;
        RECT 83.870 72.840 84.040 73.010 ;
        RECT 84.230 72.840 84.400 73.010 ;
        RECT 84.590 72.840 84.760 73.010 ;
        RECT 84.950 72.840 85.120 73.010 ;
        RECT 85.310 72.840 85.480 73.010 ;
        RECT 85.670 72.840 85.840 73.010 ;
        RECT 86.030 72.840 86.200 73.010 ;
        RECT 86.390 72.840 86.560 73.010 ;
        RECT 86.900 72.840 87.070 73.010 ;
        RECT 87.260 72.840 87.430 73.010 ;
        RECT 87.620 72.840 87.790 73.010 ;
        RECT 87.980 72.840 88.150 73.010 ;
        RECT 88.340 72.840 88.510 73.010 ;
        RECT 88.700 72.840 88.870 73.010 ;
        RECT 89.060 72.840 89.230 73.010 ;
        RECT 89.420 72.840 89.590 73.010 ;
        RECT 89.780 72.840 89.950 73.010 ;
        RECT 90.140 72.840 90.310 73.010 ;
        RECT 90.500 72.840 90.670 73.010 ;
        RECT 90.860 72.840 91.030 73.010 ;
        RECT 91.220 72.840 91.390 73.010 ;
        RECT 91.580 72.840 91.750 73.010 ;
        RECT 91.940 72.840 92.110 73.010 ;
        RECT 92.300 72.840 92.470 73.010 ;
        RECT 92.660 72.840 92.830 73.010 ;
        RECT 93.020 72.840 93.190 73.010 ;
        RECT 93.380 72.840 93.550 73.010 ;
        RECT 93.740 72.840 93.910 73.010 ;
        RECT 94.100 72.840 94.270 73.010 ;
        RECT 94.460 72.840 94.630 73.010 ;
        RECT 94.820 72.840 94.990 73.010 ;
        RECT 95.180 72.840 95.350 73.010 ;
        RECT 95.540 72.840 95.710 73.010 ;
        RECT 95.900 72.840 96.070 73.010 ;
        RECT 96.260 72.840 96.430 73.010 ;
        RECT 96.620 72.840 96.790 73.010 ;
        RECT 96.980 72.840 97.150 73.010 ;
        RECT 97.340 72.840 97.510 73.010 ;
        RECT 97.700 72.840 97.870 73.010 ;
        RECT 98.060 72.840 98.230 73.010 ;
        RECT 98.420 72.840 98.590 73.010 ;
        RECT 98.780 72.840 98.950 73.010 ;
        RECT 99.140 72.840 99.310 73.010 ;
        RECT 99.500 72.840 99.670 73.010 ;
        RECT 99.860 72.840 100.030 73.010 ;
        RECT 100.220 72.840 100.390 73.010 ;
        RECT 100.580 72.840 100.750 73.010 ;
        RECT 100.940 72.840 101.110 73.010 ;
        RECT 101.300 72.840 101.470 73.010 ;
        RECT 101.660 72.840 101.830 73.010 ;
        RECT 102.020 72.840 102.190 73.010 ;
        RECT 102.380 72.840 102.550 73.010 ;
        RECT 102.740 72.840 102.910 73.010 ;
        RECT 103.100 72.840 103.270 73.010 ;
        RECT 103.460 72.840 103.630 73.010 ;
        RECT 103.820 72.840 103.990 73.010 ;
        RECT 104.180 72.840 104.350 73.010 ;
        RECT 104.540 72.840 104.710 73.010 ;
        RECT 104.900 72.840 105.070 73.010 ;
        RECT 105.260 72.840 105.430 73.010 ;
        RECT 105.620 72.840 105.790 73.010 ;
        RECT 105.980 72.840 106.150 73.010 ;
        RECT 106.340 72.840 106.510 73.010 ;
        RECT 106.700 72.840 106.870 73.010 ;
        RECT 107.060 72.840 107.230 73.010 ;
        RECT 107.420 72.840 107.590 73.010 ;
        RECT 107.780 72.840 107.950 73.010 ;
        RECT 108.140 72.840 108.310 73.010 ;
        RECT 108.500 72.840 108.670 73.010 ;
        RECT 108.860 72.840 109.030 73.010 ;
        RECT 109.220 72.840 109.390 73.010 ;
        RECT 109.580 72.840 109.750 73.010 ;
        RECT 109.940 72.840 110.110 73.010 ;
        RECT 110.300 72.840 110.470 73.010 ;
        RECT 110.660 72.840 110.830 73.010 ;
        RECT 111.020 72.840 111.190 73.010 ;
        RECT 111.380 72.840 111.550 73.010 ;
        RECT 111.740 72.840 111.910 73.010 ;
        RECT 112.100 72.840 112.270 73.010 ;
        RECT 112.460 72.840 112.630 73.010 ;
        RECT 112.820 72.840 112.990 73.010 ;
        RECT 113.180 72.840 113.350 73.010 ;
        RECT 113.540 72.840 113.710 73.010 ;
        RECT 113.900 72.840 114.070 73.010 ;
        RECT 114.260 72.840 114.430 73.010 ;
        RECT 114.620 72.840 114.790 73.010 ;
        RECT 114.980 72.840 115.150 73.010 ;
        RECT 115.340 72.840 115.510 73.010 ;
        RECT 115.700 72.840 115.870 73.010 ;
        RECT 116.060 72.840 116.230 73.010 ;
        RECT 116.420 72.840 116.590 73.010 ;
        RECT 116.780 72.840 116.950 73.010 ;
        RECT 117.140 72.840 117.310 73.010 ;
        RECT 117.500 72.840 117.670 73.010 ;
        RECT 117.860 72.840 118.030 73.010 ;
        RECT 118.220 72.840 118.390 73.010 ;
        RECT 118.580 72.840 118.750 73.010 ;
        RECT 118.940 72.840 119.110 73.010 ;
        RECT 119.300 72.840 119.470 73.010 ;
        RECT 119.660 72.840 119.830 73.010 ;
        RECT 120.020 72.840 120.190 73.010 ;
        RECT 120.380 72.840 120.550 73.010 ;
        RECT 120.740 72.840 120.910 73.010 ;
        RECT 121.100 72.840 121.270 73.010 ;
        RECT 121.460 72.840 121.630 73.010 ;
        RECT 121.820 72.840 121.990 73.010 ;
        RECT 122.180 72.840 122.350 73.010 ;
        RECT 122.540 72.840 122.710 73.010 ;
        RECT 122.900 72.840 123.070 73.010 ;
        RECT 123.260 72.840 123.430 73.010 ;
        RECT 123.620 72.840 123.790 73.010 ;
        RECT 123.980 72.840 124.150 73.010 ;
        RECT 124.340 72.840 124.510 73.010 ;
        RECT 124.700 72.840 124.870 73.010 ;
        RECT 125.060 72.840 125.230 73.010 ;
        RECT 125.420 72.840 125.590 73.010 ;
        RECT 125.780 72.840 125.950 73.010 ;
        RECT 126.140 72.840 126.310 73.010 ;
        RECT 126.500 72.840 126.670 73.010 ;
        RECT 126.860 72.840 127.030 73.010 ;
        RECT 127.220 72.840 127.390 73.010 ;
        RECT 127.580 72.840 127.750 73.010 ;
        RECT 127.940 72.840 128.110 73.010 ;
        RECT 128.300 72.840 128.470 73.010 ;
        RECT 128.660 72.840 128.830 73.010 ;
        RECT 129.020 72.840 129.190 73.010 ;
        RECT 129.380 72.840 129.550 73.010 ;
        RECT 129.740 72.840 129.910 73.010 ;
        RECT 130.100 72.840 130.270 73.010 ;
        RECT 130.670 72.900 130.840 73.070 ;
        RECT 137.130 74.595 137.300 74.765 ;
        RECT 137.530 74.655 137.700 74.825 ;
        RECT 137.890 74.655 138.060 74.825 ;
        RECT 138.250 74.655 138.420 74.825 ;
        RECT 138.610 74.655 138.780 74.825 ;
        RECT 138.970 74.655 139.140 74.825 ;
        RECT 139.330 74.655 139.500 74.825 ;
        RECT 139.690 74.655 139.860 74.825 ;
        RECT 140.050 74.655 140.220 74.825 ;
        RECT 140.410 74.655 140.580 74.825 ;
        RECT 140.770 74.655 140.940 74.825 ;
        RECT 141.130 74.655 141.300 74.825 ;
        RECT 141.490 74.655 141.660 74.825 ;
        RECT 141.850 74.655 142.020 74.825 ;
        RECT 137.130 74.235 137.300 74.405 ;
        RECT 137.130 73.875 137.300 74.045 ;
        RECT 139.090 74.105 139.260 74.275 ;
        RECT 139.950 74.105 140.120 74.275 ;
        RECT 141.910 74.210 142.080 74.380 ;
        RECT 137.130 73.515 137.300 73.685 ;
        RECT 137.130 73.155 137.300 73.325 ;
        RECT 137.800 73.600 137.970 73.770 ;
        RECT 137.800 73.240 137.970 73.410 ;
        RECT 138.230 73.600 138.400 73.770 ;
        RECT 138.230 73.240 138.400 73.410 ;
        RECT 138.660 73.600 138.830 73.770 ;
        RECT 138.660 73.240 138.830 73.410 ;
        RECT 139.090 73.600 139.260 73.770 ;
        RECT 139.090 73.240 139.260 73.410 ;
        RECT 139.520 73.600 139.690 73.770 ;
        RECT 139.520 73.240 139.690 73.410 ;
        RECT 139.950 73.600 140.120 73.770 ;
        RECT 139.950 73.240 140.120 73.410 ;
        RECT 140.380 73.600 140.550 73.770 ;
        RECT 140.380 73.240 140.550 73.410 ;
        RECT 140.810 73.600 140.980 73.770 ;
        RECT 140.810 73.240 140.980 73.410 ;
        RECT 141.240 73.600 141.410 73.770 ;
        RECT 141.240 73.240 141.410 73.410 ;
        RECT 141.910 73.850 142.080 74.020 ;
        RECT 141.910 73.490 142.080 73.660 ;
        RECT 141.910 73.130 142.080 73.300 ;
        RECT 137.130 72.795 137.300 72.965 ;
        RECT 138.230 72.735 138.400 72.905 ;
        RECT 140.810 72.735 140.980 72.905 ;
        RECT 141.910 72.770 142.080 72.940 ;
        RECT 137.130 72.435 137.300 72.605 ;
        RECT 89.560 71.905 89.730 72.075 ;
        RECT 90.080 71.965 90.250 72.135 ;
        RECT 90.440 71.965 90.610 72.135 ;
        RECT 90.800 71.965 90.970 72.135 ;
        RECT 91.160 71.965 91.330 72.135 ;
        RECT 91.520 71.965 91.690 72.135 ;
        RECT 91.880 71.965 92.050 72.135 ;
        RECT 92.240 71.965 92.410 72.135 ;
        RECT 92.600 71.965 92.770 72.135 ;
        RECT 92.960 71.965 93.130 72.135 ;
        RECT 93.320 71.965 93.490 72.135 ;
        RECT 93.680 71.965 93.850 72.135 ;
        RECT 94.040 71.965 94.210 72.135 ;
        RECT 94.400 71.965 94.570 72.135 ;
        RECT 94.760 71.965 94.930 72.135 ;
        RECT 95.120 71.965 95.290 72.135 ;
        RECT 95.480 71.965 95.650 72.135 ;
        RECT 95.840 71.965 96.010 72.135 ;
        RECT 96.200 71.965 96.370 72.135 ;
        RECT 96.560 71.965 96.730 72.135 ;
        RECT 96.920 71.965 97.090 72.135 ;
        RECT 97.280 71.965 97.450 72.135 ;
        RECT 97.640 71.965 97.810 72.135 ;
        RECT 89.560 71.545 89.730 71.715 ;
        RECT 89.560 71.185 89.730 71.355 ;
        RECT 93.200 71.415 93.370 71.585 ;
        RECT 94.060 71.415 94.230 71.585 ;
        RECT 97.700 71.415 97.870 71.585 ;
        RECT 89.560 70.825 89.730 70.995 ;
        RECT 89.560 70.465 89.730 70.635 ;
        RECT 89.560 70.105 89.730 70.275 ;
        RECT 90.190 70.760 90.360 70.930 ;
        RECT 90.190 70.400 90.360 70.570 ;
        RECT 90.620 70.760 90.790 70.930 ;
        RECT 90.620 70.400 90.790 70.570 ;
        RECT 91.050 70.760 91.220 70.930 ;
        RECT 91.050 70.400 91.220 70.570 ;
        RECT 91.480 70.760 91.650 70.930 ;
        RECT 91.480 70.400 91.650 70.570 ;
        RECT 91.910 70.760 92.080 70.930 ;
        RECT 91.910 70.400 92.080 70.570 ;
        RECT 92.340 70.760 92.510 70.930 ;
        RECT 92.340 70.400 92.510 70.570 ;
        RECT 92.770 70.760 92.940 70.930 ;
        RECT 92.770 70.400 92.940 70.570 ;
        RECT 93.200 70.760 93.370 70.930 ;
        RECT 93.200 70.400 93.370 70.570 ;
        RECT 93.630 70.760 93.800 70.930 ;
        RECT 93.630 70.400 93.800 70.570 ;
        RECT 94.060 70.760 94.230 70.930 ;
        RECT 94.060 70.400 94.230 70.570 ;
        RECT 94.490 70.760 94.660 70.930 ;
        RECT 94.490 70.400 94.660 70.570 ;
        RECT 94.920 70.760 95.090 70.930 ;
        RECT 94.920 70.400 95.090 70.570 ;
        RECT 95.350 70.760 95.520 70.930 ;
        RECT 95.350 70.400 95.520 70.570 ;
        RECT 95.780 70.760 95.950 70.930 ;
        RECT 95.780 70.400 95.950 70.570 ;
        RECT 96.210 70.760 96.380 70.930 ;
        RECT 96.210 70.400 96.380 70.570 ;
        RECT 96.640 70.760 96.810 70.930 ;
        RECT 96.640 70.400 96.810 70.570 ;
        RECT 97.070 70.760 97.240 70.930 ;
        RECT 97.070 70.400 97.240 70.570 ;
        RECT 97.700 71.055 97.870 71.225 ;
        RECT 97.700 70.695 97.870 70.865 ;
        RECT 97.700 70.335 97.870 70.505 ;
        RECT 89.560 69.745 89.730 69.915 ;
        RECT 90.620 69.745 90.790 69.915 ;
        RECT 91.480 69.745 91.650 69.915 ;
        RECT 92.340 69.745 92.510 69.915 ;
        RECT 94.920 69.745 95.090 69.915 ;
        RECT 95.780 69.745 95.950 69.915 ;
        RECT 96.640 69.745 96.810 69.915 ;
        RECT 97.700 69.975 97.870 70.145 ;
        RECT 97.700 69.615 97.870 69.785 ;
        RECT 89.620 69.195 89.790 69.365 ;
        RECT 89.980 69.195 90.150 69.365 ;
        RECT 90.340 69.195 90.510 69.365 ;
        RECT 90.700 69.195 90.870 69.365 ;
        RECT 91.060 69.195 91.230 69.365 ;
        RECT 91.420 69.195 91.590 69.365 ;
        RECT 91.780 69.195 91.950 69.365 ;
        RECT 92.140 69.195 92.310 69.365 ;
        RECT 92.500 69.195 92.670 69.365 ;
        RECT 92.860 69.195 93.030 69.365 ;
        RECT 93.220 69.195 93.390 69.365 ;
        RECT 93.810 69.195 93.980 69.365 ;
        RECT 94.170 69.195 94.340 69.365 ;
        RECT 94.530 69.195 94.700 69.365 ;
        RECT 94.890 69.195 95.060 69.365 ;
        RECT 95.250 69.195 95.420 69.365 ;
        RECT 95.610 69.195 95.780 69.365 ;
        RECT 95.970 69.195 96.140 69.365 ;
        RECT 96.330 69.195 96.500 69.365 ;
        RECT 96.690 69.195 96.860 69.365 ;
        RECT 97.050 69.195 97.220 69.365 ;
        RECT 97.700 69.255 97.870 69.425 ;
        RECT 123.760 71.905 123.930 72.075 ;
        RECT 124.280 71.965 124.450 72.135 ;
        RECT 124.640 71.965 124.810 72.135 ;
        RECT 125.000 71.965 125.170 72.135 ;
        RECT 125.360 71.965 125.530 72.135 ;
        RECT 125.720 71.965 125.890 72.135 ;
        RECT 126.080 71.965 126.250 72.135 ;
        RECT 126.440 71.965 126.610 72.135 ;
        RECT 126.800 71.965 126.970 72.135 ;
        RECT 127.160 71.965 127.330 72.135 ;
        RECT 127.520 71.965 127.690 72.135 ;
        RECT 127.880 71.965 128.050 72.135 ;
        RECT 128.240 71.965 128.410 72.135 ;
        RECT 128.600 71.965 128.770 72.135 ;
        RECT 128.960 71.965 129.130 72.135 ;
        RECT 129.320 71.965 129.490 72.135 ;
        RECT 129.680 71.965 129.850 72.135 ;
        RECT 130.040 71.965 130.210 72.135 ;
        RECT 130.400 71.965 130.570 72.135 ;
        RECT 130.760 71.965 130.930 72.135 ;
        RECT 131.120 71.965 131.290 72.135 ;
        RECT 131.480 71.965 131.650 72.135 ;
        RECT 131.840 71.965 132.010 72.135 ;
        RECT 123.760 71.545 123.930 71.715 ;
        RECT 123.760 71.185 123.930 71.355 ;
        RECT 127.400 71.415 127.570 71.585 ;
        RECT 128.260 71.415 128.430 71.585 ;
        RECT 131.900 71.415 132.070 71.585 ;
        RECT 123.760 70.825 123.930 70.995 ;
        RECT 123.760 70.465 123.930 70.635 ;
        RECT 123.760 70.105 123.930 70.275 ;
        RECT 124.390 70.760 124.560 70.930 ;
        RECT 124.390 70.400 124.560 70.570 ;
        RECT 124.820 70.760 124.990 70.930 ;
        RECT 124.820 70.400 124.990 70.570 ;
        RECT 125.250 70.760 125.420 70.930 ;
        RECT 125.250 70.400 125.420 70.570 ;
        RECT 125.680 70.760 125.850 70.930 ;
        RECT 125.680 70.400 125.850 70.570 ;
        RECT 126.110 70.760 126.280 70.930 ;
        RECT 126.110 70.400 126.280 70.570 ;
        RECT 126.540 70.760 126.710 70.930 ;
        RECT 126.540 70.400 126.710 70.570 ;
        RECT 126.970 70.760 127.140 70.930 ;
        RECT 126.970 70.400 127.140 70.570 ;
        RECT 127.400 70.760 127.570 70.930 ;
        RECT 127.400 70.400 127.570 70.570 ;
        RECT 127.830 70.760 128.000 70.930 ;
        RECT 127.830 70.400 128.000 70.570 ;
        RECT 128.260 70.760 128.430 70.930 ;
        RECT 128.260 70.400 128.430 70.570 ;
        RECT 128.690 70.760 128.860 70.930 ;
        RECT 128.690 70.400 128.860 70.570 ;
        RECT 129.120 70.760 129.290 70.930 ;
        RECT 129.120 70.400 129.290 70.570 ;
        RECT 129.550 70.760 129.720 70.930 ;
        RECT 129.550 70.400 129.720 70.570 ;
        RECT 129.980 70.760 130.150 70.930 ;
        RECT 129.980 70.400 130.150 70.570 ;
        RECT 130.410 70.760 130.580 70.930 ;
        RECT 130.410 70.400 130.580 70.570 ;
        RECT 130.840 70.760 131.010 70.930 ;
        RECT 130.840 70.400 131.010 70.570 ;
        RECT 131.270 70.760 131.440 70.930 ;
        RECT 131.270 70.400 131.440 70.570 ;
        RECT 131.900 71.055 132.070 71.225 ;
        RECT 131.900 70.695 132.070 70.865 ;
        RECT 131.900 70.335 132.070 70.505 ;
        RECT 123.760 69.745 123.930 69.915 ;
        RECT 124.820 69.745 124.990 69.915 ;
        RECT 125.680 69.745 125.850 69.915 ;
        RECT 126.540 69.745 126.710 69.915 ;
        RECT 129.120 69.745 129.290 69.915 ;
        RECT 129.980 69.745 130.150 69.915 ;
        RECT 130.840 69.745 131.010 69.915 ;
        RECT 131.900 69.975 132.070 70.145 ;
        RECT 131.900 69.615 132.070 69.785 ;
        RECT 137.130 71.880 137.300 72.050 ;
        RECT 137.130 71.520 137.300 71.690 ;
        RECT 141.910 72.410 142.080 72.580 ;
        RECT 141.910 72.050 142.080 72.220 ;
        RECT 141.910 71.690 142.080 71.860 ;
        RECT 137.130 71.160 137.300 71.330 ;
        RECT 139.090 71.390 139.260 71.560 ;
        RECT 139.950 71.390 140.120 71.560 ;
        RECT 141.910 71.330 142.080 71.500 ;
        RECT 137.130 70.800 137.300 70.970 ;
        RECT 137.130 70.440 137.300 70.610 ;
        RECT 137.800 70.885 137.970 71.055 ;
        RECT 137.800 70.525 137.970 70.695 ;
        RECT 138.230 70.885 138.400 71.055 ;
        RECT 138.230 70.525 138.400 70.695 ;
        RECT 138.660 70.885 138.830 71.055 ;
        RECT 138.660 70.525 138.830 70.695 ;
        RECT 139.090 70.885 139.260 71.055 ;
        RECT 139.090 70.525 139.260 70.695 ;
        RECT 139.520 70.885 139.690 71.055 ;
        RECT 139.520 70.525 139.690 70.695 ;
        RECT 139.950 70.885 140.120 71.055 ;
        RECT 139.950 70.525 140.120 70.695 ;
        RECT 140.380 70.885 140.550 71.055 ;
        RECT 140.380 70.525 140.550 70.695 ;
        RECT 140.810 70.885 140.980 71.055 ;
        RECT 140.810 70.525 140.980 70.695 ;
        RECT 141.240 70.885 141.410 71.055 ;
        RECT 141.240 70.525 141.410 70.695 ;
        RECT 141.910 70.970 142.080 71.140 ;
        RECT 141.910 70.610 142.080 70.780 ;
        RECT 137.130 70.080 137.300 70.250 ;
        RECT 138.230 70.020 138.400 70.190 ;
        RECT 140.810 70.020 140.980 70.190 ;
        RECT 141.910 70.250 142.080 70.420 ;
        RECT 141.910 69.890 142.080 70.060 ;
        RECT 137.190 69.470 137.360 69.640 ;
        RECT 137.550 69.470 137.720 69.640 ;
        RECT 137.910 69.470 138.080 69.640 ;
        RECT 138.270 69.470 138.440 69.640 ;
        RECT 138.630 69.470 138.800 69.640 ;
        RECT 138.990 69.470 139.160 69.640 ;
        RECT 139.350 69.470 139.520 69.640 ;
        RECT 139.710 69.470 139.880 69.640 ;
        RECT 140.070 69.470 140.240 69.640 ;
        RECT 140.430 69.470 140.600 69.640 ;
        RECT 140.790 69.470 140.960 69.640 ;
        RECT 141.150 69.470 141.320 69.640 ;
        RECT 141.510 69.470 141.680 69.640 ;
        RECT 141.910 69.530 142.080 69.700 ;
        RECT 142.420 74.595 142.590 74.765 ;
        RECT 143.100 74.655 143.270 74.825 ;
        RECT 143.460 74.655 143.630 74.825 ;
        RECT 143.820 74.655 143.990 74.825 ;
        RECT 144.180 74.655 144.350 74.825 ;
        RECT 144.540 74.655 144.710 74.825 ;
        RECT 144.900 74.655 145.070 74.825 ;
        RECT 145.260 74.655 145.430 74.825 ;
        RECT 145.620 74.655 145.790 74.825 ;
        RECT 145.980 74.655 146.150 74.825 ;
        RECT 146.340 74.655 146.510 74.825 ;
        RECT 146.700 74.655 146.870 74.825 ;
        RECT 147.060 74.655 147.230 74.825 ;
        RECT 142.420 74.235 142.590 74.405 ;
        RECT 142.420 73.875 142.590 74.045 ;
        RECT 144.340 74.105 144.510 74.275 ;
        RECT 145.200 74.105 145.370 74.275 ;
        RECT 147.120 74.210 147.290 74.380 ;
        RECT 142.420 73.515 142.590 73.685 ;
        RECT 142.420 73.155 142.590 73.325 ;
        RECT 143.050 73.600 143.220 73.770 ;
        RECT 143.050 73.240 143.220 73.410 ;
        RECT 143.480 73.600 143.650 73.770 ;
        RECT 143.480 73.240 143.650 73.410 ;
        RECT 143.910 73.600 144.080 73.770 ;
        RECT 143.910 73.240 144.080 73.410 ;
        RECT 144.340 73.600 144.510 73.770 ;
        RECT 144.340 73.240 144.510 73.410 ;
        RECT 144.770 73.600 144.940 73.770 ;
        RECT 144.770 73.240 144.940 73.410 ;
        RECT 145.200 73.600 145.370 73.770 ;
        RECT 145.200 73.240 145.370 73.410 ;
        RECT 145.630 73.600 145.800 73.770 ;
        RECT 145.630 73.240 145.800 73.410 ;
        RECT 146.060 73.600 146.230 73.770 ;
        RECT 146.060 73.240 146.230 73.410 ;
        RECT 146.490 73.600 146.660 73.770 ;
        RECT 146.490 73.240 146.660 73.410 ;
        RECT 147.120 73.850 147.290 74.020 ;
        RECT 147.120 73.490 147.290 73.660 ;
        RECT 147.120 73.130 147.290 73.300 ;
        RECT 142.420 72.795 142.590 72.965 ;
        RECT 143.480 72.735 143.650 72.905 ;
        RECT 146.060 72.735 146.230 72.905 ;
        RECT 147.120 72.770 147.290 72.940 ;
        RECT 142.420 72.435 142.590 72.605 ;
        RECT 142.420 71.880 142.590 72.050 ;
        RECT 142.420 71.520 142.590 71.690 ;
        RECT 147.120 72.410 147.290 72.580 ;
        RECT 147.120 72.050 147.290 72.220 ;
        RECT 147.120 71.690 147.290 71.860 ;
        RECT 142.420 71.160 142.590 71.330 ;
        RECT 144.340 71.390 144.510 71.560 ;
        RECT 145.200 71.390 145.370 71.560 ;
        RECT 147.120 71.330 147.290 71.500 ;
        RECT 142.420 70.800 142.590 70.970 ;
        RECT 142.420 70.440 142.590 70.610 ;
        RECT 143.050 70.885 143.220 71.055 ;
        RECT 143.050 70.525 143.220 70.695 ;
        RECT 143.480 70.885 143.650 71.055 ;
        RECT 143.480 70.525 143.650 70.695 ;
        RECT 143.910 70.885 144.080 71.055 ;
        RECT 143.910 70.525 144.080 70.695 ;
        RECT 144.340 70.885 144.510 71.055 ;
        RECT 144.340 70.525 144.510 70.695 ;
        RECT 144.770 70.885 144.940 71.055 ;
        RECT 144.770 70.525 144.940 70.695 ;
        RECT 145.200 70.885 145.370 71.055 ;
        RECT 145.200 70.525 145.370 70.695 ;
        RECT 145.630 70.885 145.800 71.055 ;
        RECT 145.630 70.525 145.800 70.695 ;
        RECT 146.060 70.885 146.230 71.055 ;
        RECT 146.060 70.525 146.230 70.695 ;
        RECT 146.490 70.885 146.660 71.055 ;
        RECT 146.490 70.525 146.660 70.695 ;
        RECT 147.120 70.970 147.290 71.140 ;
        RECT 147.120 70.610 147.290 70.780 ;
        RECT 142.420 70.080 142.590 70.250 ;
        RECT 143.480 70.020 143.650 70.190 ;
        RECT 146.060 70.020 146.230 70.190 ;
        RECT 147.120 70.250 147.290 70.420 ;
        RECT 147.120 69.890 147.290 70.060 ;
        RECT 142.480 69.470 142.650 69.640 ;
        RECT 142.840 69.470 143.010 69.640 ;
        RECT 143.200 69.470 143.370 69.640 ;
        RECT 143.560 69.470 143.730 69.640 ;
        RECT 143.920 69.470 144.090 69.640 ;
        RECT 144.280 69.470 144.450 69.640 ;
        RECT 144.640 69.470 144.810 69.640 ;
        RECT 145.000 69.470 145.170 69.640 ;
        RECT 145.360 69.470 145.530 69.640 ;
        RECT 145.720 69.470 145.890 69.640 ;
        RECT 146.080 69.470 146.250 69.640 ;
        RECT 146.440 69.470 146.610 69.640 ;
        RECT 147.120 69.530 147.290 69.700 ;
        RECT 123.820 69.195 123.990 69.365 ;
        RECT 124.180 69.195 124.350 69.365 ;
        RECT 124.540 69.195 124.710 69.365 ;
        RECT 124.900 69.195 125.070 69.365 ;
        RECT 125.260 69.195 125.430 69.365 ;
        RECT 125.620 69.195 125.790 69.365 ;
        RECT 125.980 69.195 126.150 69.365 ;
        RECT 126.340 69.195 126.510 69.365 ;
        RECT 126.700 69.195 126.870 69.365 ;
        RECT 127.060 69.195 127.230 69.365 ;
        RECT 127.420 69.195 127.590 69.365 ;
        RECT 128.010 69.195 128.180 69.365 ;
        RECT 128.370 69.195 128.540 69.365 ;
        RECT 128.730 69.195 128.900 69.365 ;
        RECT 129.090 69.195 129.260 69.365 ;
        RECT 129.450 69.195 129.620 69.365 ;
        RECT 129.810 69.195 129.980 69.365 ;
        RECT 130.170 69.195 130.340 69.365 ;
        RECT 130.530 69.195 130.700 69.365 ;
        RECT 130.890 69.195 131.060 69.365 ;
        RECT 131.250 69.195 131.420 69.365 ;
        RECT 131.900 69.255 132.070 69.425 ;
        RECT 89.325 68.335 89.495 68.505 ;
        RECT 89.865 68.395 90.035 68.565 ;
        RECT 90.225 68.395 90.395 68.565 ;
        RECT 90.585 68.395 90.755 68.565 ;
        RECT 90.945 68.395 91.115 68.565 ;
        RECT 91.305 68.395 91.475 68.565 ;
        RECT 91.665 68.395 91.835 68.565 ;
        RECT 92.025 68.395 92.195 68.565 ;
        RECT 92.385 68.395 92.555 68.565 ;
        RECT 92.745 68.395 92.915 68.565 ;
        RECT 93.105 68.395 93.275 68.565 ;
        RECT 89.325 67.975 89.495 68.145 ;
        RECT 89.325 67.615 89.495 67.785 ;
        RECT 90.385 67.845 90.555 68.015 ;
        RECT 92.105 67.845 92.275 68.015 ;
        RECT 93.165 67.785 93.335 67.955 ;
        RECT 89.325 67.255 89.495 67.425 ;
        RECT 89.325 66.895 89.495 67.065 ;
        RECT 89.955 67.340 90.125 67.510 ;
        RECT 89.955 66.980 90.125 67.150 ;
        RECT 90.385 67.340 90.555 67.510 ;
        RECT 90.385 66.980 90.555 67.150 ;
        RECT 90.815 67.340 90.985 67.510 ;
        RECT 90.815 66.980 90.985 67.150 ;
        RECT 91.245 67.340 91.415 67.510 ;
        RECT 91.245 66.980 91.415 67.150 ;
        RECT 91.675 67.340 91.845 67.510 ;
        RECT 91.675 66.980 91.845 67.150 ;
        RECT 92.105 67.340 92.275 67.510 ;
        RECT 92.105 66.980 92.275 67.150 ;
        RECT 92.535 67.340 92.705 67.510 ;
        RECT 92.535 66.980 92.705 67.150 ;
        RECT 93.165 67.425 93.335 67.595 ;
        RECT 93.165 67.065 93.335 67.235 ;
        RECT 89.325 66.535 89.495 66.705 ;
        RECT 91.245 66.475 91.415 66.645 ;
        RECT 93.165 66.705 93.335 66.875 ;
        RECT 93.165 66.345 93.335 66.515 ;
        RECT 89.385 65.925 89.555 66.095 ;
        RECT 89.745 65.925 89.915 66.095 ;
        RECT 90.105 65.925 90.275 66.095 ;
        RECT 90.465 65.925 90.635 66.095 ;
        RECT 90.825 65.925 90.995 66.095 ;
        RECT 91.425 65.925 91.595 66.095 ;
        RECT 91.785 65.925 91.955 66.095 ;
        RECT 92.145 65.925 92.315 66.095 ;
        RECT 92.505 65.925 92.675 66.095 ;
        RECT 93.165 65.985 93.335 66.155 ;
        RECT 93.955 68.335 94.125 68.505 ;
        RECT 94.575 68.395 94.745 68.565 ;
        RECT 94.935 68.395 95.105 68.565 ;
        RECT 95.295 68.395 95.465 68.565 ;
        RECT 95.655 68.395 95.825 68.565 ;
        RECT 96.015 68.395 96.185 68.565 ;
        RECT 96.375 68.395 96.545 68.565 ;
        RECT 96.735 68.395 96.905 68.565 ;
        RECT 97.095 68.395 97.265 68.565 ;
        RECT 97.455 68.395 97.625 68.565 ;
        RECT 97.815 68.395 97.985 68.565 ;
        RECT 93.955 67.975 94.125 68.145 ;
        RECT 93.955 67.615 94.125 67.785 ;
        RECT 95.915 67.845 96.085 68.015 ;
        RECT 97.875 67.785 98.045 67.955 ;
        RECT 93.955 67.255 94.125 67.425 ;
        RECT 93.955 66.895 94.125 67.065 ;
        RECT 94.625 67.340 94.795 67.510 ;
        RECT 94.625 66.980 94.795 67.150 ;
        RECT 95.055 67.340 95.225 67.510 ;
        RECT 95.055 66.980 95.225 67.150 ;
        RECT 95.485 67.340 95.655 67.510 ;
        RECT 95.485 66.980 95.655 67.150 ;
        RECT 95.915 67.340 96.085 67.510 ;
        RECT 95.915 66.980 96.085 67.150 ;
        RECT 96.345 67.340 96.515 67.510 ;
        RECT 96.345 66.980 96.515 67.150 ;
        RECT 96.775 67.340 96.945 67.510 ;
        RECT 96.775 66.980 96.945 67.150 ;
        RECT 97.205 67.340 97.375 67.510 ;
        RECT 97.205 66.980 97.375 67.150 ;
        RECT 97.875 67.425 98.045 67.595 ;
        RECT 97.875 67.065 98.045 67.235 ;
        RECT 93.955 66.535 94.125 66.705 ;
        RECT 95.055 66.475 95.225 66.645 ;
        RECT 96.775 66.475 96.945 66.645 ;
        RECT 97.875 66.705 98.045 66.875 ;
        RECT 97.875 66.345 98.045 66.515 ;
        RECT 94.015 65.925 94.185 66.095 ;
        RECT 94.375 65.925 94.545 66.095 ;
        RECT 94.735 65.925 94.905 66.095 ;
        RECT 95.095 65.925 95.265 66.095 ;
        RECT 95.455 65.925 95.625 66.095 ;
        RECT 96.095 65.925 96.265 66.095 ;
        RECT 96.455 65.925 96.625 66.095 ;
        RECT 96.815 65.925 96.985 66.095 ;
        RECT 97.175 65.925 97.345 66.095 ;
        RECT 97.875 65.985 98.045 66.155 ;
        RECT 123.525 68.335 123.695 68.505 ;
        RECT 124.065 68.395 124.235 68.565 ;
        RECT 124.425 68.395 124.595 68.565 ;
        RECT 124.785 68.395 124.955 68.565 ;
        RECT 125.145 68.395 125.315 68.565 ;
        RECT 125.505 68.395 125.675 68.565 ;
        RECT 125.865 68.395 126.035 68.565 ;
        RECT 126.225 68.395 126.395 68.565 ;
        RECT 126.585 68.395 126.755 68.565 ;
        RECT 126.945 68.395 127.115 68.565 ;
        RECT 127.305 68.395 127.475 68.565 ;
        RECT 123.525 67.975 123.695 68.145 ;
        RECT 123.525 67.615 123.695 67.785 ;
        RECT 124.585 67.845 124.755 68.015 ;
        RECT 126.305 67.845 126.475 68.015 ;
        RECT 127.365 67.785 127.535 67.955 ;
        RECT 123.525 67.255 123.695 67.425 ;
        RECT 123.525 66.895 123.695 67.065 ;
        RECT 124.155 67.340 124.325 67.510 ;
        RECT 124.155 66.980 124.325 67.150 ;
        RECT 124.585 67.340 124.755 67.510 ;
        RECT 124.585 66.980 124.755 67.150 ;
        RECT 125.015 67.340 125.185 67.510 ;
        RECT 125.015 66.980 125.185 67.150 ;
        RECT 125.445 67.340 125.615 67.510 ;
        RECT 125.445 66.980 125.615 67.150 ;
        RECT 125.875 67.340 126.045 67.510 ;
        RECT 125.875 66.980 126.045 67.150 ;
        RECT 126.305 67.340 126.475 67.510 ;
        RECT 126.305 66.980 126.475 67.150 ;
        RECT 126.735 67.340 126.905 67.510 ;
        RECT 126.735 66.980 126.905 67.150 ;
        RECT 127.365 67.425 127.535 67.595 ;
        RECT 127.365 67.065 127.535 67.235 ;
        RECT 123.525 66.535 123.695 66.705 ;
        RECT 125.445 66.475 125.615 66.645 ;
        RECT 127.365 66.705 127.535 66.875 ;
        RECT 127.365 66.345 127.535 66.515 ;
        RECT 123.585 65.925 123.755 66.095 ;
        RECT 123.945 65.925 124.115 66.095 ;
        RECT 124.305 65.925 124.475 66.095 ;
        RECT 124.665 65.925 124.835 66.095 ;
        RECT 125.025 65.925 125.195 66.095 ;
        RECT 125.625 65.925 125.795 66.095 ;
        RECT 125.985 65.925 126.155 66.095 ;
        RECT 126.345 65.925 126.515 66.095 ;
        RECT 126.705 65.925 126.875 66.095 ;
        RECT 127.365 65.985 127.535 66.155 ;
        RECT 128.155 68.335 128.325 68.505 ;
        RECT 128.775 68.395 128.945 68.565 ;
        RECT 129.135 68.395 129.305 68.565 ;
        RECT 129.495 68.395 129.665 68.565 ;
        RECT 129.855 68.395 130.025 68.565 ;
        RECT 130.215 68.395 130.385 68.565 ;
        RECT 130.575 68.395 130.745 68.565 ;
        RECT 130.935 68.395 131.105 68.565 ;
        RECT 131.295 68.395 131.465 68.565 ;
        RECT 131.655 68.395 131.825 68.565 ;
        RECT 132.015 68.395 132.185 68.565 ;
        RECT 128.155 67.975 128.325 68.145 ;
        RECT 128.155 67.615 128.325 67.785 ;
        RECT 130.115 67.845 130.285 68.015 ;
        RECT 132.075 67.785 132.245 67.955 ;
        RECT 128.155 67.255 128.325 67.425 ;
        RECT 128.155 66.895 128.325 67.065 ;
        RECT 128.825 67.340 128.995 67.510 ;
        RECT 128.825 66.980 128.995 67.150 ;
        RECT 129.255 67.340 129.425 67.510 ;
        RECT 129.255 66.980 129.425 67.150 ;
        RECT 129.685 67.340 129.855 67.510 ;
        RECT 129.685 66.980 129.855 67.150 ;
        RECT 130.115 67.340 130.285 67.510 ;
        RECT 130.115 66.980 130.285 67.150 ;
        RECT 130.545 67.340 130.715 67.510 ;
        RECT 130.545 66.980 130.715 67.150 ;
        RECT 130.975 67.340 131.145 67.510 ;
        RECT 130.975 66.980 131.145 67.150 ;
        RECT 131.405 67.340 131.575 67.510 ;
        RECT 131.405 66.980 131.575 67.150 ;
        RECT 132.075 67.425 132.245 67.595 ;
        RECT 132.075 67.065 132.245 67.235 ;
        RECT 128.155 66.535 128.325 66.705 ;
        RECT 129.255 66.475 129.425 66.645 ;
        RECT 130.975 66.475 131.145 66.645 ;
        RECT 132.075 66.705 132.245 66.875 ;
        RECT 132.075 66.345 132.245 66.515 ;
        RECT 128.215 65.925 128.385 66.095 ;
        RECT 128.575 65.925 128.745 66.095 ;
        RECT 128.935 65.925 129.105 66.095 ;
        RECT 129.295 65.925 129.465 66.095 ;
        RECT 129.655 65.925 129.825 66.095 ;
        RECT 130.295 65.925 130.465 66.095 ;
        RECT 130.655 65.925 130.825 66.095 ;
        RECT 131.015 65.925 131.185 66.095 ;
        RECT 131.375 65.925 131.545 66.095 ;
        RECT 132.075 65.985 132.245 66.155 ;
        RECT 136.850 68.185 137.020 68.355 ;
        RECT 137.530 68.245 137.700 68.415 ;
        RECT 137.890 68.245 138.060 68.415 ;
        RECT 138.250 68.245 138.420 68.415 ;
        RECT 138.610 68.245 138.780 68.415 ;
        RECT 138.970 68.245 139.140 68.415 ;
        RECT 139.330 68.245 139.500 68.415 ;
        RECT 139.690 68.245 139.860 68.415 ;
        RECT 140.050 68.245 140.220 68.415 ;
        RECT 140.410 68.245 140.580 68.415 ;
        RECT 140.770 68.245 140.940 68.415 ;
        RECT 141.130 68.245 141.300 68.415 ;
        RECT 141.490 68.245 141.660 68.415 ;
        RECT 141.850 68.245 142.020 68.415 ;
        RECT 142.210 68.245 142.380 68.415 ;
        RECT 142.570 68.245 142.740 68.415 ;
        RECT 142.930 68.245 143.100 68.415 ;
        RECT 143.290 68.245 143.460 68.415 ;
        RECT 143.650 68.245 143.820 68.415 ;
        RECT 144.010 68.245 144.180 68.415 ;
        RECT 144.370 68.245 144.540 68.415 ;
        RECT 144.730 68.245 144.900 68.415 ;
        RECT 145.090 68.245 145.260 68.415 ;
        RECT 145.450 68.245 145.620 68.415 ;
        RECT 145.810 68.245 145.980 68.415 ;
        RECT 146.170 68.245 146.340 68.415 ;
        RECT 146.530 68.245 146.700 68.415 ;
        RECT 146.890 68.245 147.060 68.415 ;
        RECT 147.250 68.245 147.420 68.415 ;
        RECT 136.850 67.825 137.020 67.995 ;
        RECT 136.850 67.465 137.020 67.635 ;
        RECT 137.940 67.695 138.110 67.865 ;
        RECT 138.300 67.695 138.470 67.865 ;
        RECT 138.660 67.695 138.830 67.865 ;
        RECT 139.020 67.695 139.190 67.865 ;
        RECT 139.380 67.695 139.550 67.865 ;
        RECT 144.780 67.695 144.950 67.865 ;
        RECT 145.140 67.695 145.310 67.865 ;
        RECT 145.500 67.695 145.670 67.865 ;
        RECT 145.860 67.695 146.030 67.865 ;
        RECT 146.220 67.695 146.390 67.865 ;
        RECT 147.310 67.635 147.480 67.805 ;
        RECT 136.850 67.105 137.020 67.275 ;
        RECT 136.850 66.745 137.020 66.915 ;
        RECT 137.520 67.190 137.690 67.360 ;
        RECT 137.520 66.830 137.690 67.000 ;
        RECT 139.800 67.190 139.970 67.360 ;
        RECT 139.800 66.830 139.970 67.000 ;
        RECT 142.080 67.190 142.250 67.360 ;
        RECT 142.080 66.830 142.250 67.000 ;
        RECT 144.360 67.190 144.530 67.360 ;
        RECT 144.360 66.830 144.530 67.000 ;
        RECT 146.640 67.190 146.810 67.360 ;
        RECT 146.640 66.830 146.810 67.000 ;
        RECT 147.310 67.275 147.480 67.445 ;
        RECT 147.310 66.915 147.480 67.085 ;
        RECT 136.850 66.385 137.020 66.555 ;
        RECT 140.220 66.325 140.390 66.495 ;
        RECT 140.580 66.325 140.750 66.495 ;
        RECT 140.940 66.325 141.110 66.495 ;
        RECT 141.300 66.325 141.470 66.495 ;
        RECT 141.660 66.325 141.830 66.495 ;
        RECT 142.500 66.325 142.670 66.495 ;
        RECT 142.860 66.325 143.030 66.495 ;
        RECT 143.220 66.325 143.390 66.495 ;
        RECT 143.580 66.325 143.750 66.495 ;
        RECT 143.940 66.325 144.110 66.495 ;
        RECT 147.310 66.555 147.480 66.725 ;
        RECT 147.310 66.195 147.480 66.365 ;
        RECT 136.910 65.775 137.080 65.945 ;
        RECT 137.270 65.775 137.440 65.945 ;
        RECT 137.630 65.775 137.800 65.945 ;
        RECT 137.990 65.775 138.160 65.945 ;
        RECT 138.350 65.775 138.520 65.945 ;
        RECT 138.710 65.775 138.880 65.945 ;
        RECT 139.070 65.775 139.240 65.945 ;
        RECT 139.430 65.775 139.600 65.945 ;
        RECT 139.790 65.775 139.960 65.945 ;
        RECT 140.150 65.775 140.320 65.945 ;
        RECT 140.510 65.775 140.680 65.945 ;
        RECT 140.870 65.775 141.040 65.945 ;
        RECT 141.230 65.775 141.400 65.945 ;
        RECT 141.590 65.775 141.760 65.945 ;
        RECT 142.260 65.775 142.430 65.945 ;
        RECT 142.620 65.775 142.790 65.945 ;
        RECT 142.980 65.775 143.150 65.945 ;
        RECT 143.340 65.775 143.510 65.945 ;
        RECT 143.700 65.775 143.870 65.945 ;
        RECT 144.060 65.775 144.230 65.945 ;
        RECT 144.420 65.775 144.590 65.945 ;
        RECT 144.780 65.775 144.950 65.945 ;
        RECT 145.140 65.775 145.310 65.945 ;
        RECT 145.500 65.775 145.670 65.945 ;
        RECT 145.860 65.775 146.030 65.945 ;
        RECT 146.220 65.775 146.390 65.945 ;
        RECT 146.580 65.775 146.750 65.945 ;
        RECT 146.940 65.775 147.110 65.945 ;
        RECT 147.310 65.835 147.480 66.005 ;
        RECT 33.930 65.005 34.100 65.175 ;
        RECT 34.290 65.005 34.460 65.175 ;
        RECT 34.650 65.005 34.820 65.175 ;
        RECT 35.010 65.005 35.180 65.175 ;
        RECT 35.370 65.005 35.540 65.175 ;
        RECT 35.730 65.005 35.900 65.175 ;
        RECT 36.090 65.005 36.260 65.175 ;
        RECT 36.450 65.005 36.620 65.175 ;
        RECT 36.810 65.005 36.980 65.175 ;
        RECT 37.170 65.005 37.340 65.175 ;
        RECT 37.530 65.005 37.700 65.175 ;
        RECT 37.890 65.005 38.060 65.175 ;
        RECT 33.580 64.705 33.750 64.875 ;
        RECT 38.360 64.705 38.530 64.875 ;
        RECT 33.580 64.345 33.750 64.515 ;
        RECT 33.580 63.985 33.750 64.155 ;
        RECT 33.580 63.625 33.750 63.795 ;
        RECT 33.580 63.265 33.750 63.435 ;
        RECT 33.580 62.905 33.750 63.075 ;
        RECT 33.580 62.545 33.750 62.715 ;
        RECT 34.250 64.180 34.420 64.350 ;
        RECT 34.250 63.820 34.420 63.990 ;
        RECT 34.250 63.460 34.420 63.630 ;
        RECT 34.250 63.100 34.420 63.270 ;
        RECT 34.250 62.740 34.420 62.910 ;
        RECT 34.680 64.180 34.850 64.350 ;
        RECT 34.680 63.820 34.850 63.990 ;
        RECT 34.680 63.460 34.850 63.630 ;
        RECT 34.680 63.100 34.850 63.270 ;
        RECT 34.680 62.740 34.850 62.910 ;
        RECT 35.110 64.180 35.280 64.350 ;
        RECT 35.110 63.820 35.280 63.990 ;
        RECT 35.110 63.460 35.280 63.630 ;
        RECT 35.110 63.100 35.280 63.270 ;
        RECT 35.110 62.740 35.280 62.910 ;
        RECT 35.540 64.180 35.710 64.350 ;
        RECT 35.540 63.820 35.710 63.990 ;
        RECT 35.540 63.460 35.710 63.630 ;
        RECT 35.540 63.100 35.710 63.270 ;
        RECT 35.540 62.740 35.710 62.910 ;
        RECT 35.970 64.180 36.140 64.350 ;
        RECT 35.970 63.820 36.140 63.990 ;
        RECT 35.970 63.460 36.140 63.630 ;
        RECT 35.970 63.100 36.140 63.270 ;
        RECT 35.970 62.740 36.140 62.910 ;
        RECT 36.400 64.180 36.570 64.350 ;
        RECT 36.400 63.820 36.570 63.990 ;
        RECT 36.400 63.460 36.570 63.630 ;
        RECT 36.400 63.100 36.570 63.270 ;
        RECT 36.400 62.740 36.570 62.910 ;
        RECT 36.830 64.180 37.000 64.350 ;
        RECT 36.830 63.820 37.000 63.990 ;
        RECT 36.830 63.460 37.000 63.630 ;
        RECT 36.830 63.100 37.000 63.270 ;
        RECT 36.830 62.740 37.000 62.910 ;
        RECT 37.260 64.180 37.430 64.350 ;
        RECT 37.260 63.820 37.430 63.990 ;
        RECT 37.260 63.460 37.430 63.630 ;
        RECT 37.260 63.100 37.430 63.270 ;
        RECT 37.260 62.740 37.430 62.910 ;
        RECT 37.690 64.180 37.860 64.350 ;
        RECT 37.690 63.820 37.860 63.990 ;
        RECT 37.690 63.460 37.860 63.630 ;
        RECT 37.690 63.100 37.860 63.270 ;
        RECT 37.690 62.740 37.860 62.910 ;
        RECT 38.360 64.345 38.530 64.515 ;
        RECT 38.360 63.985 38.530 64.155 ;
        RECT 38.360 63.625 38.530 63.795 ;
        RECT 38.360 63.265 38.530 63.435 ;
        RECT 38.360 62.905 38.530 63.075 ;
        RECT 38.360 62.545 38.530 62.715 ;
        RECT 33.580 62.185 33.750 62.355 ;
        RECT 34.500 62.125 34.670 62.295 ;
        RECT 34.860 62.125 35.030 62.295 ;
        RECT 35.360 62.125 35.530 62.295 ;
        RECT 35.720 62.125 35.890 62.295 ;
        RECT 36.220 62.125 36.390 62.295 ;
        RECT 36.580 62.125 36.750 62.295 ;
        RECT 37.080 62.125 37.250 62.295 ;
        RECT 37.440 62.125 37.610 62.295 ;
        RECT 38.360 62.185 38.530 62.355 ;
        RECT 42.730 64.785 42.900 64.955 ;
        RECT 43.170 64.845 43.340 65.015 ;
        RECT 43.530 64.845 43.700 65.015 ;
        RECT 43.890 64.845 44.060 65.015 ;
        RECT 44.250 64.845 44.420 65.015 ;
        RECT 44.610 64.845 44.780 65.015 ;
        RECT 44.970 64.845 45.140 65.015 ;
        RECT 45.330 64.845 45.500 65.015 ;
        RECT 45.690 64.845 45.860 65.015 ;
        RECT 46.050 64.845 46.220 65.015 ;
        RECT 46.410 64.845 46.580 65.015 ;
        RECT 46.770 64.845 46.940 65.015 ;
        RECT 47.130 64.845 47.300 65.015 ;
        RECT 47.490 64.845 47.660 65.015 ;
        RECT 47.850 64.845 48.020 65.015 ;
        RECT 48.210 64.845 48.380 65.015 ;
        RECT 48.570 64.845 48.740 65.015 ;
        RECT 48.930 64.845 49.100 65.015 ;
        RECT 49.290 64.845 49.460 65.015 ;
        RECT 49.650 64.845 49.820 65.015 ;
        RECT 50.010 64.845 50.180 65.015 ;
        RECT 50.370 64.845 50.540 65.015 ;
        RECT 50.730 64.845 50.900 65.015 ;
        RECT 51.090 64.845 51.260 65.015 ;
        RECT 51.450 64.845 51.620 65.015 ;
        RECT 51.810 64.845 51.980 65.015 ;
        RECT 52.170 64.845 52.340 65.015 ;
        RECT 52.530 64.845 52.700 65.015 ;
        RECT 52.890 64.845 53.060 65.015 ;
        RECT 53.250 64.845 53.420 65.015 ;
        RECT 53.610 64.845 53.780 65.015 ;
        RECT 53.970 64.845 54.140 65.015 ;
        RECT 54.330 64.845 54.500 65.015 ;
        RECT 54.690 64.845 54.860 65.015 ;
        RECT 55.050 64.845 55.220 65.015 ;
        RECT 55.410 64.845 55.580 65.015 ;
        RECT 55.770 64.845 55.940 65.015 ;
        RECT 56.130 64.845 56.300 65.015 ;
        RECT 56.490 64.845 56.660 65.015 ;
        RECT 56.850 64.845 57.020 65.015 ;
        RECT 57.210 64.845 57.380 65.015 ;
        RECT 57.570 64.845 57.740 65.015 ;
        RECT 57.930 64.845 58.100 65.015 ;
        RECT 58.290 64.845 58.460 65.015 ;
        RECT 58.650 64.845 58.820 65.015 ;
        RECT 59.010 64.845 59.180 65.015 ;
        RECT 59.370 64.845 59.540 65.015 ;
        RECT 59.730 64.845 59.900 65.015 ;
        RECT 60.090 64.845 60.260 65.015 ;
        RECT 60.450 64.845 60.620 65.015 ;
        RECT 60.810 64.845 60.980 65.015 ;
        RECT 61.170 64.845 61.340 65.015 ;
        RECT 61.530 64.845 61.700 65.015 ;
        RECT 61.890 64.845 62.060 65.015 ;
        RECT 62.250 64.845 62.420 65.015 ;
        RECT 62.610 64.845 62.780 65.015 ;
        RECT 62.970 64.845 63.140 65.015 ;
        RECT 63.330 64.845 63.500 65.015 ;
        RECT 63.690 64.845 63.860 65.015 ;
        RECT 64.050 64.845 64.220 65.015 ;
        RECT 64.410 64.845 64.580 65.015 ;
        RECT 64.770 64.845 64.940 65.015 ;
        RECT 65.130 64.845 65.300 65.015 ;
        RECT 65.490 64.845 65.660 65.015 ;
        RECT 65.850 64.845 66.020 65.015 ;
        RECT 66.210 64.845 66.380 65.015 ;
        RECT 66.570 64.845 66.740 65.015 ;
        RECT 66.930 64.845 67.100 65.015 ;
        RECT 67.290 64.845 67.460 65.015 ;
        RECT 67.650 64.845 67.820 65.015 ;
        RECT 68.010 64.845 68.180 65.015 ;
        RECT 68.370 64.845 68.540 65.015 ;
        RECT 68.730 64.845 68.900 65.015 ;
        RECT 69.090 64.845 69.260 65.015 ;
        RECT 69.450 64.845 69.620 65.015 ;
        RECT 69.810 64.845 69.980 65.015 ;
        RECT 70.170 64.845 70.340 65.015 ;
        RECT 70.530 64.845 70.700 65.015 ;
        RECT 70.890 64.845 71.060 65.015 ;
        RECT 71.250 64.845 71.420 65.015 ;
        RECT 71.610 64.845 71.780 65.015 ;
        RECT 71.970 64.845 72.140 65.015 ;
        RECT 72.330 64.845 72.500 65.015 ;
        RECT 72.690 64.845 72.860 65.015 ;
        RECT 73.050 64.845 73.220 65.015 ;
        RECT 73.410 64.845 73.580 65.015 ;
        RECT 73.770 64.845 73.940 65.015 ;
        RECT 74.130 64.845 74.300 65.015 ;
        RECT 74.490 64.845 74.660 65.015 ;
        RECT 74.850 64.845 75.020 65.015 ;
        RECT 75.210 64.845 75.380 65.015 ;
        RECT 75.570 64.845 75.740 65.015 ;
        RECT 75.930 64.845 76.100 65.015 ;
        RECT 76.290 64.845 76.460 65.015 ;
        RECT 76.650 64.845 76.820 65.015 ;
        RECT 77.010 64.845 77.180 65.015 ;
        RECT 77.370 64.845 77.540 65.015 ;
        RECT 77.730 64.845 77.900 65.015 ;
        RECT 78.090 64.845 78.260 65.015 ;
        RECT 78.450 64.845 78.620 65.015 ;
        RECT 78.810 64.845 78.980 65.015 ;
        RECT 79.170 64.845 79.340 65.015 ;
        RECT 79.530 64.845 79.700 65.015 ;
        RECT 79.890 64.845 80.060 65.015 ;
        RECT 80.250 64.845 80.420 65.015 ;
        RECT 80.610 64.845 80.780 65.015 ;
        RECT 80.970 64.845 81.140 65.015 ;
        RECT 81.330 64.845 81.500 65.015 ;
        RECT 81.690 64.845 81.860 65.015 ;
        RECT 82.050 64.845 82.220 65.015 ;
        RECT 82.410 64.845 82.580 65.015 ;
        RECT 82.770 64.845 82.940 65.015 ;
        RECT 83.130 64.845 83.300 65.015 ;
        RECT 83.490 64.845 83.660 65.015 ;
        RECT 83.850 64.845 84.020 65.015 ;
        RECT 84.210 64.845 84.380 65.015 ;
        RECT 84.570 64.845 84.740 65.015 ;
        RECT 84.930 64.845 85.100 65.015 ;
        RECT 85.290 64.845 85.460 65.015 ;
        RECT 85.650 64.845 85.820 65.015 ;
        RECT 86.010 64.845 86.180 65.015 ;
        RECT 86.370 64.845 86.540 65.015 ;
        RECT 86.730 64.845 86.900 65.015 ;
        RECT 87.090 64.845 87.260 65.015 ;
        RECT 87.450 64.845 87.620 65.015 ;
        RECT 87.810 64.845 87.980 65.015 ;
        RECT 88.170 64.845 88.340 65.015 ;
        RECT 88.530 64.845 88.700 65.015 ;
        RECT 88.890 64.845 89.060 65.015 ;
        RECT 89.250 64.845 89.420 65.015 ;
        RECT 89.610 64.845 89.780 65.015 ;
        RECT 89.970 64.845 90.140 65.015 ;
        RECT 90.330 64.845 90.500 65.015 ;
        RECT 90.690 64.845 90.860 65.015 ;
        RECT 91.050 64.845 91.220 65.015 ;
        RECT 91.410 64.845 91.580 65.015 ;
        RECT 91.770 64.845 91.940 65.015 ;
        RECT 92.130 64.845 92.300 65.015 ;
        RECT 92.490 64.845 92.660 65.015 ;
        RECT 92.850 64.845 93.020 65.015 ;
        RECT 93.210 64.845 93.380 65.015 ;
        RECT 93.570 64.845 93.740 65.015 ;
        RECT 93.930 64.845 94.100 65.015 ;
        RECT 94.290 64.845 94.460 65.015 ;
        RECT 94.650 64.845 94.820 65.015 ;
        RECT 95.010 64.845 95.180 65.015 ;
        RECT 95.370 64.845 95.540 65.015 ;
        RECT 95.730 64.845 95.900 65.015 ;
        RECT 96.090 64.845 96.260 65.015 ;
        RECT 96.450 64.845 96.620 65.015 ;
        RECT 96.810 64.845 96.980 65.015 ;
        RECT 97.170 64.845 97.340 65.015 ;
        RECT 97.530 64.845 97.700 65.015 ;
        RECT 97.890 64.845 98.060 65.015 ;
        RECT 98.250 64.845 98.420 65.015 ;
        RECT 98.610 64.845 98.780 65.015 ;
        RECT 98.970 64.845 99.140 65.015 ;
        RECT 99.330 64.845 99.500 65.015 ;
        RECT 99.690 64.845 99.860 65.015 ;
        RECT 100.050 64.845 100.220 65.015 ;
        RECT 100.410 64.845 100.580 65.015 ;
        RECT 100.770 64.845 100.940 65.015 ;
        RECT 101.130 64.845 101.300 65.015 ;
        RECT 101.490 64.845 101.660 65.015 ;
        RECT 101.850 64.845 102.020 65.015 ;
        RECT 102.210 64.845 102.380 65.015 ;
        RECT 102.570 64.845 102.740 65.015 ;
        RECT 102.930 64.845 103.100 65.015 ;
        RECT 103.290 64.845 103.460 65.015 ;
        RECT 103.650 64.845 103.820 65.015 ;
        RECT 104.010 64.845 104.180 65.015 ;
        RECT 104.370 64.845 104.540 65.015 ;
        RECT 104.730 64.845 104.900 65.015 ;
        RECT 105.090 64.845 105.260 65.015 ;
        RECT 105.450 64.845 105.620 65.015 ;
        RECT 105.810 64.845 105.980 65.015 ;
        RECT 106.170 64.845 106.340 65.015 ;
        RECT 106.530 64.845 106.700 65.015 ;
        RECT 106.890 64.845 107.060 65.015 ;
        RECT 107.250 64.845 107.420 65.015 ;
        RECT 107.610 64.845 107.780 65.015 ;
        RECT 107.970 64.845 108.140 65.015 ;
        RECT 108.330 64.845 108.500 65.015 ;
        RECT 108.690 64.845 108.860 65.015 ;
        RECT 109.050 64.845 109.220 65.015 ;
        RECT 109.410 64.845 109.580 65.015 ;
        RECT 109.770 64.845 109.940 65.015 ;
        RECT 110.130 64.845 110.300 65.015 ;
        RECT 110.490 64.845 110.660 65.015 ;
        RECT 110.850 64.845 111.020 65.015 ;
        RECT 111.210 64.845 111.380 65.015 ;
        RECT 111.570 64.845 111.740 65.015 ;
        RECT 111.930 64.845 112.100 65.015 ;
        RECT 112.290 64.845 112.460 65.015 ;
        RECT 112.650 64.845 112.820 65.015 ;
        RECT 113.010 64.845 113.180 65.015 ;
        RECT 113.370 64.845 113.540 65.015 ;
        RECT 113.730 64.845 113.900 65.015 ;
        RECT 114.090 64.845 114.260 65.015 ;
        RECT 114.450 64.845 114.620 65.015 ;
        RECT 114.810 64.845 114.980 65.015 ;
        RECT 115.170 64.845 115.340 65.015 ;
        RECT 115.530 64.845 115.700 65.015 ;
        RECT 115.890 64.845 116.060 65.015 ;
        RECT 116.250 64.845 116.420 65.015 ;
        RECT 116.610 64.845 116.780 65.015 ;
        RECT 116.970 64.845 117.140 65.015 ;
        RECT 117.330 64.845 117.500 65.015 ;
        RECT 117.690 64.845 117.860 65.015 ;
        RECT 118.050 64.845 118.220 65.015 ;
        RECT 118.410 64.845 118.580 65.015 ;
        RECT 118.770 64.845 118.940 65.015 ;
        RECT 119.130 64.845 119.300 65.015 ;
        RECT 119.490 64.845 119.660 65.015 ;
        RECT 119.850 64.845 120.020 65.015 ;
        RECT 120.210 64.845 120.380 65.015 ;
        RECT 120.570 64.845 120.740 65.015 ;
        RECT 120.930 64.845 121.100 65.015 ;
        RECT 121.290 64.845 121.460 65.015 ;
        RECT 121.650 64.845 121.820 65.015 ;
        RECT 122.010 64.845 122.180 65.015 ;
        RECT 122.370 64.845 122.540 65.015 ;
        RECT 122.730 64.845 122.900 65.015 ;
        RECT 123.090 64.845 123.260 65.015 ;
        RECT 123.450 64.845 123.620 65.015 ;
        RECT 123.810 64.845 123.980 65.015 ;
        RECT 124.170 64.845 124.340 65.015 ;
        RECT 124.530 64.845 124.700 65.015 ;
        RECT 124.890 64.845 125.060 65.015 ;
        RECT 125.250 64.845 125.420 65.015 ;
        RECT 125.610 64.845 125.780 65.015 ;
        RECT 125.970 64.845 126.140 65.015 ;
        RECT 126.330 64.845 126.500 65.015 ;
        RECT 126.690 64.845 126.860 65.015 ;
        RECT 127.050 64.845 127.220 65.015 ;
        RECT 127.410 64.845 127.580 65.015 ;
        RECT 127.770 64.845 127.940 65.015 ;
        RECT 128.130 64.845 128.300 65.015 ;
        RECT 128.490 64.845 128.660 65.015 ;
        RECT 128.850 64.845 129.020 65.015 ;
        RECT 129.210 64.845 129.380 65.015 ;
        RECT 129.570 64.845 129.740 65.015 ;
        RECT 129.930 64.845 130.100 65.015 ;
        RECT 130.290 64.845 130.460 65.015 ;
        RECT 130.650 64.845 130.820 65.015 ;
        RECT 131.010 64.845 131.180 65.015 ;
        RECT 131.370 64.845 131.540 65.015 ;
        RECT 131.730 64.845 131.900 65.015 ;
        RECT 132.090 64.845 132.260 65.015 ;
        RECT 132.450 64.845 132.620 65.015 ;
        RECT 132.810 64.845 132.980 65.015 ;
        RECT 133.170 64.845 133.340 65.015 ;
        RECT 133.530 64.845 133.700 65.015 ;
        RECT 133.890 64.845 134.060 65.015 ;
        RECT 134.250 64.845 134.420 65.015 ;
        RECT 134.610 64.845 134.780 65.015 ;
        RECT 134.970 64.845 135.140 65.015 ;
        RECT 135.330 64.845 135.500 65.015 ;
        RECT 135.690 64.845 135.860 65.015 ;
        RECT 136.050 64.845 136.220 65.015 ;
        RECT 136.410 64.845 136.580 65.015 ;
        RECT 136.770 64.845 136.940 65.015 ;
        RECT 137.130 64.845 137.300 65.015 ;
        RECT 137.490 64.845 137.660 65.015 ;
        RECT 137.850 64.845 138.020 65.015 ;
        RECT 138.210 64.845 138.380 65.015 ;
        RECT 138.570 64.845 138.740 65.015 ;
        RECT 138.930 64.845 139.100 65.015 ;
        RECT 139.290 64.845 139.460 65.015 ;
        RECT 139.650 64.845 139.820 65.015 ;
        RECT 140.010 64.845 140.180 65.015 ;
        RECT 140.370 64.845 140.540 65.015 ;
        RECT 140.730 64.845 140.900 65.015 ;
        RECT 141.090 64.845 141.260 65.015 ;
        RECT 141.450 64.845 141.620 65.015 ;
        RECT 141.810 64.845 141.980 65.015 ;
        RECT 142.170 64.845 142.340 65.015 ;
        RECT 142.530 64.845 142.700 65.015 ;
        RECT 142.890 64.845 143.060 65.015 ;
        RECT 143.250 64.845 143.420 65.015 ;
        RECT 143.610 64.845 143.780 65.015 ;
        RECT 143.970 64.845 144.140 65.015 ;
        RECT 144.330 64.845 144.500 65.015 ;
        RECT 42.730 64.425 42.900 64.595 ;
        RECT 42.730 64.065 42.900 64.235 ;
        RECT 144.390 64.375 144.560 64.545 ;
        RECT 42.730 63.705 42.900 63.875 ;
        RECT 42.730 63.345 42.900 63.515 ;
        RECT 43.400 63.790 43.570 63.960 ;
        RECT 43.400 63.430 43.570 63.600 ;
        RECT 45.680 63.790 45.850 63.960 ;
        RECT 45.680 63.430 45.850 63.600 ;
        RECT 47.960 63.790 48.130 63.960 ;
        RECT 47.960 63.430 48.130 63.600 ;
        RECT 50.240 63.790 50.410 63.960 ;
        RECT 50.240 63.430 50.410 63.600 ;
        RECT 52.520 63.790 52.690 63.960 ;
        RECT 52.520 63.430 52.690 63.600 ;
        RECT 54.800 63.790 54.970 63.960 ;
        RECT 54.800 63.430 54.970 63.600 ;
        RECT 57.080 63.790 57.250 63.960 ;
        RECT 57.080 63.430 57.250 63.600 ;
        RECT 59.360 63.790 59.530 63.960 ;
        RECT 59.360 63.430 59.530 63.600 ;
        RECT 61.640 63.790 61.810 63.960 ;
        RECT 61.640 63.430 61.810 63.600 ;
        RECT 63.920 63.790 64.090 63.960 ;
        RECT 63.920 63.430 64.090 63.600 ;
        RECT 66.200 63.790 66.370 63.960 ;
        RECT 66.200 63.430 66.370 63.600 ;
        RECT 68.480 63.790 68.650 63.960 ;
        RECT 68.480 63.430 68.650 63.600 ;
        RECT 70.760 63.790 70.930 63.960 ;
        RECT 70.760 63.430 70.930 63.600 ;
        RECT 73.040 63.790 73.210 63.960 ;
        RECT 73.040 63.430 73.210 63.600 ;
        RECT 75.320 63.790 75.490 63.960 ;
        RECT 75.320 63.430 75.490 63.600 ;
        RECT 77.600 63.790 77.770 63.960 ;
        RECT 77.600 63.430 77.770 63.600 ;
        RECT 79.880 63.790 80.050 63.960 ;
        RECT 79.880 63.430 80.050 63.600 ;
        RECT 82.160 63.790 82.330 63.960 ;
        RECT 82.160 63.430 82.330 63.600 ;
        RECT 84.440 63.790 84.610 63.960 ;
        RECT 84.440 63.430 84.610 63.600 ;
        RECT 86.720 63.790 86.890 63.960 ;
        RECT 86.720 63.430 86.890 63.600 ;
        RECT 89.000 63.790 89.170 63.960 ;
        RECT 89.000 63.430 89.170 63.600 ;
        RECT 91.280 63.790 91.450 63.960 ;
        RECT 91.280 63.430 91.450 63.600 ;
        RECT 93.560 63.790 93.730 63.960 ;
        RECT 93.560 63.430 93.730 63.600 ;
        RECT 95.840 63.790 96.010 63.960 ;
        RECT 95.840 63.430 96.010 63.600 ;
        RECT 98.120 63.790 98.290 63.960 ;
        RECT 98.120 63.430 98.290 63.600 ;
        RECT 100.400 63.790 100.570 63.960 ;
        RECT 100.400 63.430 100.570 63.600 ;
        RECT 102.680 63.790 102.850 63.960 ;
        RECT 102.680 63.430 102.850 63.600 ;
        RECT 104.960 63.790 105.130 63.960 ;
        RECT 104.960 63.430 105.130 63.600 ;
        RECT 107.240 63.790 107.410 63.960 ;
        RECT 107.240 63.430 107.410 63.600 ;
        RECT 109.520 63.790 109.690 63.960 ;
        RECT 109.520 63.430 109.690 63.600 ;
        RECT 111.800 63.790 111.970 63.960 ;
        RECT 111.800 63.430 111.970 63.600 ;
        RECT 114.080 63.790 114.250 63.960 ;
        RECT 114.080 63.430 114.250 63.600 ;
        RECT 116.360 63.790 116.530 63.960 ;
        RECT 116.360 63.430 116.530 63.600 ;
        RECT 118.640 63.790 118.810 63.960 ;
        RECT 118.640 63.430 118.810 63.600 ;
        RECT 120.920 63.790 121.090 63.960 ;
        RECT 120.920 63.430 121.090 63.600 ;
        RECT 123.200 63.790 123.370 63.960 ;
        RECT 123.200 63.430 123.370 63.600 ;
        RECT 125.480 63.790 125.650 63.960 ;
        RECT 125.480 63.430 125.650 63.600 ;
        RECT 127.760 63.790 127.930 63.960 ;
        RECT 127.760 63.430 127.930 63.600 ;
        RECT 130.040 63.790 130.210 63.960 ;
        RECT 130.040 63.430 130.210 63.600 ;
        RECT 132.320 63.790 132.490 63.960 ;
        RECT 132.320 63.430 132.490 63.600 ;
        RECT 134.600 63.790 134.770 63.960 ;
        RECT 134.600 63.430 134.770 63.600 ;
        RECT 136.880 63.790 137.050 63.960 ;
        RECT 136.880 63.430 137.050 63.600 ;
        RECT 139.160 63.790 139.330 63.960 ;
        RECT 139.160 63.430 139.330 63.600 ;
        RECT 141.440 63.790 141.610 63.960 ;
        RECT 141.440 63.430 141.610 63.600 ;
        RECT 143.720 63.790 143.890 63.960 ;
        RECT 143.720 63.430 143.890 63.600 ;
        RECT 144.390 64.015 144.560 64.185 ;
        RECT 144.390 63.655 144.560 63.825 ;
        RECT 144.390 63.295 144.560 63.465 ;
        RECT 42.730 62.985 42.900 63.155 ;
        RECT 43.820 62.925 43.990 63.095 ;
        RECT 44.180 62.925 44.350 63.095 ;
        RECT 44.540 62.925 44.710 63.095 ;
        RECT 44.900 62.925 45.070 63.095 ;
        RECT 45.260 62.925 45.430 63.095 ;
        RECT 46.100 62.925 46.270 63.095 ;
        RECT 46.460 62.925 46.630 63.095 ;
        RECT 46.820 62.925 46.990 63.095 ;
        RECT 47.180 62.925 47.350 63.095 ;
        RECT 47.540 62.925 47.710 63.095 ;
        RECT 48.380 62.925 48.550 63.095 ;
        RECT 48.740 62.925 48.910 63.095 ;
        RECT 49.100 62.925 49.270 63.095 ;
        RECT 49.460 62.925 49.630 63.095 ;
        RECT 49.820 62.925 49.990 63.095 ;
        RECT 50.660 62.925 50.830 63.095 ;
        RECT 51.020 62.925 51.190 63.095 ;
        RECT 51.380 62.925 51.550 63.095 ;
        RECT 51.740 62.925 51.910 63.095 ;
        RECT 52.100 62.925 52.270 63.095 ;
        RECT 52.940 62.925 53.110 63.095 ;
        RECT 53.300 62.925 53.470 63.095 ;
        RECT 53.660 62.925 53.830 63.095 ;
        RECT 54.020 62.925 54.190 63.095 ;
        RECT 54.380 62.925 54.550 63.095 ;
        RECT 55.220 62.925 55.390 63.095 ;
        RECT 55.580 62.925 55.750 63.095 ;
        RECT 55.940 62.925 56.110 63.095 ;
        RECT 56.300 62.925 56.470 63.095 ;
        RECT 56.660 62.925 56.830 63.095 ;
        RECT 57.500 62.925 57.670 63.095 ;
        RECT 57.860 62.925 58.030 63.095 ;
        RECT 58.220 62.925 58.390 63.095 ;
        RECT 58.580 62.925 58.750 63.095 ;
        RECT 58.940 62.925 59.110 63.095 ;
        RECT 59.780 62.925 59.950 63.095 ;
        RECT 60.140 62.925 60.310 63.095 ;
        RECT 60.500 62.925 60.670 63.095 ;
        RECT 60.860 62.925 61.030 63.095 ;
        RECT 61.220 62.925 61.390 63.095 ;
        RECT 62.060 62.925 62.230 63.095 ;
        RECT 62.420 62.925 62.590 63.095 ;
        RECT 62.780 62.925 62.950 63.095 ;
        RECT 63.140 62.925 63.310 63.095 ;
        RECT 63.500 62.925 63.670 63.095 ;
        RECT 64.340 62.925 64.510 63.095 ;
        RECT 64.700 62.925 64.870 63.095 ;
        RECT 65.060 62.925 65.230 63.095 ;
        RECT 65.420 62.925 65.590 63.095 ;
        RECT 65.780 62.925 65.950 63.095 ;
        RECT 66.620 62.925 66.790 63.095 ;
        RECT 66.980 62.925 67.150 63.095 ;
        RECT 67.340 62.925 67.510 63.095 ;
        RECT 67.700 62.925 67.870 63.095 ;
        RECT 68.060 62.925 68.230 63.095 ;
        RECT 68.900 62.925 69.070 63.095 ;
        RECT 69.260 62.925 69.430 63.095 ;
        RECT 69.620 62.925 69.790 63.095 ;
        RECT 69.980 62.925 70.150 63.095 ;
        RECT 70.340 62.925 70.510 63.095 ;
        RECT 71.180 62.925 71.350 63.095 ;
        RECT 71.540 62.925 71.710 63.095 ;
        RECT 71.900 62.925 72.070 63.095 ;
        RECT 72.260 62.925 72.430 63.095 ;
        RECT 72.620 62.925 72.790 63.095 ;
        RECT 73.460 62.925 73.630 63.095 ;
        RECT 73.820 62.925 73.990 63.095 ;
        RECT 74.180 62.925 74.350 63.095 ;
        RECT 74.540 62.925 74.710 63.095 ;
        RECT 74.900 62.925 75.070 63.095 ;
        RECT 75.740 62.925 75.910 63.095 ;
        RECT 76.100 62.925 76.270 63.095 ;
        RECT 76.460 62.925 76.630 63.095 ;
        RECT 76.820 62.925 76.990 63.095 ;
        RECT 77.180 62.925 77.350 63.095 ;
        RECT 78.020 62.925 78.190 63.095 ;
        RECT 78.380 62.925 78.550 63.095 ;
        RECT 78.740 62.925 78.910 63.095 ;
        RECT 79.100 62.925 79.270 63.095 ;
        RECT 79.460 62.925 79.630 63.095 ;
        RECT 80.300 62.925 80.470 63.095 ;
        RECT 80.660 62.925 80.830 63.095 ;
        RECT 81.020 62.925 81.190 63.095 ;
        RECT 81.380 62.925 81.550 63.095 ;
        RECT 81.740 62.925 81.910 63.095 ;
        RECT 82.580 62.925 82.750 63.095 ;
        RECT 82.940 62.925 83.110 63.095 ;
        RECT 83.300 62.925 83.470 63.095 ;
        RECT 83.660 62.925 83.830 63.095 ;
        RECT 84.020 62.925 84.190 63.095 ;
        RECT 84.860 62.925 85.030 63.095 ;
        RECT 85.220 62.925 85.390 63.095 ;
        RECT 85.580 62.925 85.750 63.095 ;
        RECT 85.940 62.925 86.110 63.095 ;
        RECT 86.300 62.925 86.470 63.095 ;
        RECT 87.140 62.925 87.310 63.095 ;
        RECT 87.500 62.925 87.670 63.095 ;
        RECT 87.860 62.925 88.030 63.095 ;
        RECT 88.220 62.925 88.390 63.095 ;
        RECT 88.580 62.925 88.750 63.095 ;
        RECT 89.420 62.925 89.590 63.095 ;
        RECT 89.780 62.925 89.950 63.095 ;
        RECT 90.140 62.925 90.310 63.095 ;
        RECT 90.500 62.925 90.670 63.095 ;
        RECT 90.860 62.925 91.030 63.095 ;
        RECT 91.700 62.925 91.870 63.095 ;
        RECT 92.060 62.925 92.230 63.095 ;
        RECT 92.420 62.925 92.590 63.095 ;
        RECT 92.780 62.925 92.950 63.095 ;
        RECT 93.140 62.925 93.310 63.095 ;
        RECT 93.980 62.925 94.150 63.095 ;
        RECT 94.340 62.925 94.510 63.095 ;
        RECT 94.700 62.925 94.870 63.095 ;
        RECT 95.060 62.925 95.230 63.095 ;
        RECT 95.420 62.925 95.590 63.095 ;
        RECT 96.260 62.925 96.430 63.095 ;
        RECT 96.620 62.925 96.790 63.095 ;
        RECT 96.980 62.925 97.150 63.095 ;
        RECT 97.340 62.925 97.510 63.095 ;
        RECT 97.700 62.925 97.870 63.095 ;
        RECT 98.540 62.925 98.710 63.095 ;
        RECT 98.900 62.925 99.070 63.095 ;
        RECT 99.260 62.925 99.430 63.095 ;
        RECT 99.620 62.925 99.790 63.095 ;
        RECT 99.980 62.925 100.150 63.095 ;
        RECT 100.820 62.925 100.990 63.095 ;
        RECT 101.180 62.925 101.350 63.095 ;
        RECT 101.540 62.925 101.710 63.095 ;
        RECT 101.900 62.925 102.070 63.095 ;
        RECT 102.260 62.925 102.430 63.095 ;
        RECT 103.100 62.925 103.270 63.095 ;
        RECT 103.460 62.925 103.630 63.095 ;
        RECT 103.820 62.925 103.990 63.095 ;
        RECT 104.180 62.925 104.350 63.095 ;
        RECT 104.540 62.925 104.710 63.095 ;
        RECT 105.380 62.925 105.550 63.095 ;
        RECT 105.740 62.925 105.910 63.095 ;
        RECT 106.100 62.925 106.270 63.095 ;
        RECT 106.460 62.925 106.630 63.095 ;
        RECT 106.820 62.925 106.990 63.095 ;
        RECT 107.660 62.925 107.830 63.095 ;
        RECT 108.020 62.925 108.190 63.095 ;
        RECT 108.380 62.925 108.550 63.095 ;
        RECT 108.740 62.925 108.910 63.095 ;
        RECT 109.100 62.925 109.270 63.095 ;
        RECT 109.940 62.925 110.110 63.095 ;
        RECT 110.300 62.925 110.470 63.095 ;
        RECT 110.660 62.925 110.830 63.095 ;
        RECT 111.020 62.925 111.190 63.095 ;
        RECT 111.380 62.925 111.550 63.095 ;
        RECT 112.220 62.925 112.390 63.095 ;
        RECT 112.580 62.925 112.750 63.095 ;
        RECT 112.940 62.925 113.110 63.095 ;
        RECT 113.300 62.925 113.470 63.095 ;
        RECT 113.660 62.925 113.830 63.095 ;
        RECT 114.500 62.925 114.670 63.095 ;
        RECT 114.860 62.925 115.030 63.095 ;
        RECT 115.220 62.925 115.390 63.095 ;
        RECT 115.580 62.925 115.750 63.095 ;
        RECT 115.940 62.925 116.110 63.095 ;
        RECT 116.780 62.925 116.950 63.095 ;
        RECT 117.140 62.925 117.310 63.095 ;
        RECT 117.500 62.925 117.670 63.095 ;
        RECT 117.860 62.925 118.030 63.095 ;
        RECT 118.220 62.925 118.390 63.095 ;
        RECT 119.060 62.925 119.230 63.095 ;
        RECT 119.420 62.925 119.590 63.095 ;
        RECT 119.780 62.925 119.950 63.095 ;
        RECT 120.140 62.925 120.310 63.095 ;
        RECT 120.500 62.925 120.670 63.095 ;
        RECT 121.340 62.925 121.510 63.095 ;
        RECT 121.700 62.925 121.870 63.095 ;
        RECT 122.060 62.925 122.230 63.095 ;
        RECT 122.420 62.925 122.590 63.095 ;
        RECT 122.780 62.925 122.950 63.095 ;
        RECT 123.620 62.925 123.790 63.095 ;
        RECT 123.980 62.925 124.150 63.095 ;
        RECT 124.340 62.925 124.510 63.095 ;
        RECT 124.700 62.925 124.870 63.095 ;
        RECT 125.060 62.925 125.230 63.095 ;
        RECT 125.900 62.925 126.070 63.095 ;
        RECT 126.260 62.925 126.430 63.095 ;
        RECT 126.620 62.925 126.790 63.095 ;
        RECT 126.980 62.925 127.150 63.095 ;
        RECT 127.340 62.925 127.510 63.095 ;
        RECT 128.180 62.925 128.350 63.095 ;
        RECT 128.540 62.925 128.710 63.095 ;
        RECT 128.900 62.925 129.070 63.095 ;
        RECT 129.260 62.925 129.430 63.095 ;
        RECT 129.620 62.925 129.790 63.095 ;
        RECT 130.460 62.925 130.630 63.095 ;
        RECT 130.820 62.925 130.990 63.095 ;
        RECT 131.180 62.925 131.350 63.095 ;
        RECT 131.540 62.925 131.710 63.095 ;
        RECT 131.900 62.925 132.070 63.095 ;
        RECT 132.740 62.925 132.910 63.095 ;
        RECT 133.100 62.925 133.270 63.095 ;
        RECT 133.460 62.925 133.630 63.095 ;
        RECT 133.820 62.925 133.990 63.095 ;
        RECT 134.180 62.925 134.350 63.095 ;
        RECT 135.020 62.925 135.190 63.095 ;
        RECT 135.380 62.925 135.550 63.095 ;
        RECT 135.740 62.925 135.910 63.095 ;
        RECT 136.100 62.925 136.270 63.095 ;
        RECT 136.460 62.925 136.630 63.095 ;
        RECT 137.300 62.925 137.470 63.095 ;
        RECT 137.660 62.925 137.830 63.095 ;
        RECT 138.020 62.925 138.190 63.095 ;
        RECT 138.380 62.925 138.550 63.095 ;
        RECT 138.740 62.925 138.910 63.095 ;
        RECT 139.580 62.925 139.750 63.095 ;
        RECT 139.940 62.925 140.110 63.095 ;
        RECT 140.300 62.925 140.470 63.095 ;
        RECT 140.660 62.925 140.830 63.095 ;
        RECT 141.020 62.925 141.190 63.095 ;
        RECT 141.860 62.925 142.030 63.095 ;
        RECT 142.220 62.925 142.390 63.095 ;
        RECT 142.580 62.925 142.750 63.095 ;
        RECT 142.940 62.925 143.110 63.095 ;
        RECT 143.300 62.925 143.470 63.095 ;
        RECT 144.390 62.935 144.560 63.105 ;
        RECT 42.730 62.625 42.900 62.795 ;
        RECT 42.730 62.265 42.900 62.435 ;
        RECT 42.730 61.905 42.900 62.075 ;
        RECT 43.400 62.420 43.570 62.590 ;
        RECT 43.400 62.060 43.570 62.230 ;
        RECT 45.680 62.420 45.850 62.590 ;
        RECT 45.680 62.060 45.850 62.230 ;
        RECT 47.960 62.420 48.130 62.590 ;
        RECT 47.960 62.060 48.130 62.230 ;
        RECT 50.240 62.420 50.410 62.590 ;
        RECT 50.240 62.060 50.410 62.230 ;
        RECT 52.520 62.420 52.690 62.590 ;
        RECT 52.520 62.060 52.690 62.230 ;
        RECT 54.800 62.420 54.970 62.590 ;
        RECT 54.800 62.060 54.970 62.230 ;
        RECT 57.080 62.420 57.250 62.590 ;
        RECT 57.080 62.060 57.250 62.230 ;
        RECT 59.360 62.420 59.530 62.590 ;
        RECT 59.360 62.060 59.530 62.230 ;
        RECT 61.640 62.420 61.810 62.590 ;
        RECT 61.640 62.060 61.810 62.230 ;
        RECT 63.920 62.420 64.090 62.590 ;
        RECT 63.920 62.060 64.090 62.230 ;
        RECT 66.200 62.420 66.370 62.590 ;
        RECT 66.200 62.060 66.370 62.230 ;
        RECT 68.480 62.420 68.650 62.590 ;
        RECT 68.480 62.060 68.650 62.230 ;
        RECT 70.760 62.420 70.930 62.590 ;
        RECT 70.760 62.060 70.930 62.230 ;
        RECT 73.040 62.420 73.210 62.590 ;
        RECT 73.040 62.060 73.210 62.230 ;
        RECT 75.320 62.420 75.490 62.590 ;
        RECT 75.320 62.060 75.490 62.230 ;
        RECT 77.600 62.420 77.770 62.590 ;
        RECT 77.600 62.060 77.770 62.230 ;
        RECT 79.880 62.420 80.050 62.590 ;
        RECT 79.880 62.060 80.050 62.230 ;
        RECT 82.160 62.420 82.330 62.590 ;
        RECT 82.160 62.060 82.330 62.230 ;
        RECT 84.440 62.420 84.610 62.590 ;
        RECT 84.440 62.060 84.610 62.230 ;
        RECT 86.720 62.420 86.890 62.590 ;
        RECT 86.720 62.060 86.890 62.230 ;
        RECT 89.000 62.420 89.170 62.590 ;
        RECT 89.000 62.060 89.170 62.230 ;
        RECT 91.280 62.420 91.450 62.590 ;
        RECT 91.280 62.060 91.450 62.230 ;
        RECT 93.560 62.420 93.730 62.590 ;
        RECT 93.560 62.060 93.730 62.230 ;
        RECT 95.840 62.420 96.010 62.590 ;
        RECT 95.840 62.060 96.010 62.230 ;
        RECT 98.120 62.420 98.290 62.590 ;
        RECT 98.120 62.060 98.290 62.230 ;
        RECT 100.400 62.420 100.570 62.590 ;
        RECT 100.400 62.060 100.570 62.230 ;
        RECT 102.680 62.420 102.850 62.590 ;
        RECT 102.680 62.060 102.850 62.230 ;
        RECT 104.960 62.420 105.130 62.590 ;
        RECT 104.960 62.060 105.130 62.230 ;
        RECT 107.240 62.420 107.410 62.590 ;
        RECT 107.240 62.060 107.410 62.230 ;
        RECT 109.520 62.420 109.690 62.590 ;
        RECT 109.520 62.060 109.690 62.230 ;
        RECT 111.800 62.420 111.970 62.590 ;
        RECT 111.800 62.060 111.970 62.230 ;
        RECT 114.080 62.420 114.250 62.590 ;
        RECT 114.080 62.060 114.250 62.230 ;
        RECT 116.360 62.420 116.530 62.590 ;
        RECT 116.360 62.060 116.530 62.230 ;
        RECT 118.640 62.420 118.810 62.590 ;
        RECT 118.640 62.060 118.810 62.230 ;
        RECT 120.920 62.420 121.090 62.590 ;
        RECT 120.920 62.060 121.090 62.230 ;
        RECT 123.200 62.420 123.370 62.590 ;
        RECT 123.200 62.060 123.370 62.230 ;
        RECT 125.480 62.420 125.650 62.590 ;
        RECT 125.480 62.060 125.650 62.230 ;
        RECT 127.760 62.420 127.930 62.590 ;
        RECT 127.760 62.060 127.930 62.230 ;
        RECT 130.040 62.420 130.210 62.590 ;
        RECT 130.040 62.060 130.210 62.230 ;
        RECT 132.320 62.420 132.490 62.590 ;
        RECT 132.320 62.060 132.490 62.230 ;
        RECT 134.600 62.420 134.770 62.590 ;
        RECT 134.600 62.060 134.770 62.230 ;
        RECT 136.880 62.420 137.050 62.590 ;
        RECT 136.880 62.060 137.050 62.230 ;
        RECT 139.160 62.420 139.330 62.590 ;
        RECT 139.160 62.060 139.330 62.230 ;
        RECT 141.440 62.420 141.610 62.590 ;
        RECT 141.440 62.060 141.610 62.230 ;
        RECT 143.720 62.420 143.890 62.590 ;
        RECT 143.720 62.060 143.890 62.230 ;
        RECT 144.390 62.575 144.560 62.745 ;
        RECT 144.390 62.215 144.560 62.385 ;
        RECT 144.390 61.855 144.560 62.025 ;
        RECT 42.730 61.545 42.900 61.715 ;
        RECT 43.820 61.555 43.990 61.725 ;
        RECT 44.180 61.555 44.350 61.725 ;
        RECT 44.540 61.555 44.710 61.725 ;
        RECT 44.900 61.555 45.070 61.725 ;
        RECT 45.260 61.555 45.430 61.725 ;
        RECT 46.100 61.555 46.270 61.725 ;
        RECT 46.460 61.555 46.630 61.725 ;
        RECT 46.820 61.555 46.990 61.725 ;
        RECT 47.180 61.555 47.350 61.725 ;
        RECT 47.540 61.555 47.710 61.725 ;
        RECT 48.380 61.555 48.550 61.725 ;
        RECT 48.740 61.555 48.910 61.725 ;
        RECT 49.100 61.555 49.270 61.725 ;
        RECT 49.460 61.555 49.630 61.725 ;
        RECT 49.820 61.555 49.990 61.725 ;
        RECT 50.660 61.555 50.830 61.725 ;
        RECT 51.020 61.555 51.190 61.725 ;
        RECT 51.380 61.555 51.550 61.725 ;
        RECT 51.740 61.555 51.910 61.725 ;
        RECT 52.100 61.555 52.270 61.725 ;
        RECT 52.940 61.555 53.110 61.725 ;
        RECT 53.300 61.555 53.470 61.725 ;
        RECT 53.660 61.555 53.830 61.725 ;
        RECT 54.020 61.555 54.190 61.725 ;
        RECT 54.380 61.555 54.550 61.725 ;
        RECT 55.220 61.555 55.390 61.725 ;
        RECT 55.580 61.555 55.750 61.725 ;
        RECT 55.940 61.555 56.110 61.725 ;
        RECT 56.300 61.555 56.470 61.725 ;
        RECT 56.660 61.555 56.830 61.725 ;
        RECT 57.500 61.555 57.670 61.725 ;
        RECT 57.860 61.555 58.030 61.725 ;
        RECT 58.220 61.555 58.390 61.725 ;
        RECT 58.580 61.555 58.750 61.725 ;
        RECT 58.940 61.555 59.110 61.725 ;
        RECT 59.780 61.555 59.950 61.725 ;
        RECT 60.140 61.555 60.310 61.725 ;
        RECT 60.500 61.555 60.670 61.725 ;
        RECT 60.860 61.555 61.030 61.725 ;
        RECT 61.220 61.555 61.390 61.725 ;
        RECT 62.060 61.555 62.230 61.725 ;
        RECT 62.420 61.555 62.590 61.725 ;
        RECT 62.780 61.555 62.950 61.725 ;
        RECT 63.140 61.555 63.310 61.725 ;
        RECT 63.500 61.555 63.670 61.725 ;
        RECT 64.340 61.555 64.510 61.725 ;
        RECT 64.700 61.555 64.870 61.725 ;
        RECT 65.060 61.555 65.230 61.725 ;
        RECT 65.420 61.555 65.590 61.725 ;
        RECT 65.780 61.555 65.950 61.725 ;
        RECT 66.620 61.555 66.790 61.725 ;
        RECT 66.980 61.555 67.150 61.725 ;
        RECT 67.340 61.555 67.510 61.725 ;
        RECT 67.700 61.555 67.870 61.725 ;
        RECT 68.060 61.555 68.230 61.725 ;
        RECT 68.900 61.555 69.070 61.725 ;
        RECT 69.260 61.555 69.430 61.725 ;
        RECT 69.620 61.555 69.790 61.725 ;
        RECT 69.980 61.555 70.150 61.725 ;
        RECT 70.340 61.555 70.510 61.725 ;
        RECT 71.180 61.555 71.350 61.725 ;
        RECT 71.540 61.555 71.710 61.725 ;
        RECT 71.900 61.555 72.070 61.725 ;
        RECT 72.260 61.555 72.430 61.725 ;
        RECT 72.620 61.555 72.790 61.725 ;
        RECT 73.460 61.555 73.630 61.725 ;
        RECT 73.820 61.555 73.990 61.725 ;
        RECT 74.180 61.555 74.350 61.725 ;
        RECT 74.540 61.555 74.710 61.725 ;
        RECT 74.900 61.555 75.070 61.725 ;
        RECT 75.740 61.555 75.910 61.725 ;
        RECT 76.100 61.555 76.270 61.725 ;
        RECT 76.460 61.555 76.630 61.725 ;
        RECT 76.820 61.555 76.990 61.725 ;
        RECT 77.180 61.555 77.350 61.725 ;
        RECT 78.020 61.555 78.190 61.725 ;
        RECT 78.380 61.555 78.550 61.725 ;
        RECT 78.740 61.555 78.910 61.725 ;
        RECT 79.100 61.555 79.270 61.725 ;
        RECT 79.460 61.555 79.630 61.725 ;
        RECT 80.300 61.555 80.470 61.725 ;
        RECT 80.660 61.555 80.830 61.725 ;
        RECT 81.020 61.555 81.190 61.725 ;
        RECT 81.380 61.555 81.550 61.725 ;
        RECT 81.740 61.555 81.910 61.725 ;
        RECT 82.580 61.555 82.750 61.725 ;
        RECT 82.940 61.555 83.110 61.725 ;
        RECT 83.300 61.555 83.470 61.725 ;
        RECT 83.660 61.555 83.830 61.725 ;
        RECT 84.020 61.555 84.190 61.725 ;
        RECT 84.860 61.555 85.030 61.725 ;
        RECT 85.220 61.555 85.390 61.725 ;
        RECT 85.580 61.555 85.750 61.725 ;
        RECT 85.940 61.555 86.110 61.725 ;
        RECT 86.300 61.555 86.470 61.725 ;
        RECT 87.140 61.555 87.310 61.725 ;
        RECT 87.500 61.555 87.670 61.725 ;
        RECT 87.860 61.555 88.030 61.725 ;
        RECT 88.220 61.555 88.390 61.725 ;
        RECT 88.580 61.555 88.750 61.725 ;
        RECT 89.420 61.555 89.590 61.725 ;
        RECT 89.780 61.555 89.950 61.725 ;
        RECT 90.140 61.555 90.310 61.725 ;
        RECT 90.500 61.555 90.670 61.725 ;
        RECT 90.860 61.555 91.030 61.725 ;
        RECT 91.700 61.555 91.870 61.725 ;
        RECT 92.060 61.555 92.230 61.725 ;
        RECT 92.420 61.555 92.590 61.725 ;
        RECT 92.780 61.555 92.950 61.725 ;
        RECT 93.140 61.555 93.310 61.725 ;
        RECT 93.980 61.555 94.150 61.725 ;
        RECT 94.340 61.555 94.510 61.725 ;
        RECT 94.700 61.555 94.870 61.725 ;
        RECT 95.060 61.555 95.230 61.725 ;
        RECT 95.420 61.555 95.590 61.725 ;
        RECT 96.260 61.555 96.430 61.725 ;
        RECT 96.620 61.555 96.790 61.725 ;
        RECT 96.980 61.555 97.150 61.725 ;
        RECT 97.340 61.555 97.510 61.725 ;
        RECT 97.700 61.555 97.870 61.725 ;
        RECT 98.540 61.555 98.710 61.725 ;
        RECT 98.900 61.555 99.070 61.725 ;
        RECT 99.260 61.555 99.430 61.725 ;
        RECT 99.620 61.555 99.790 61.725 ;
        RECT 99.980 61.555 100.150 61.725 ;
        RECT 100.820 61.555 100.990 61.725 ;
        RECT 101.180 61.555 101.350 61.725 ;
        RECT 101.540 61.555 101.710 61.725 ;
        RECT 101.900 61.555 102.070 61.725 ;
        RECT 102.260 61.555 102.430 61.725 ;
        RECT 103.100 61.555 103.270 61.725 ;
        RECT 103.460 61.555 103.630 61.725 ;
        RECT 103.820 61.555 103.990 61.725 ;
        RECT 104.180 61.555 104.350 61.725 ;
        RECT 104.540 61.555 104.710 61.725 ;
        RECT 105.380 61.555 105.550 61.725 ;
        RECT 105.740 61.555 105.910 61.725 ;
        RECT 106.100 61.555 106.270 61.725 ;
        RECT 106.460 61.555 106.630 61.725 ;
        RECT 106.820 61.555 106.990 61.725 ;
        RECT 107.660 61.555 107.830 61.725 ;
        RECT 108.020 61.555 108.190 61.725 ;
        RECT 108.380 61.555 108.550 61.725 ;
        RECT 108.740 61.555 108.910 61.725 ;
        RECT 109.100 61.555 109.270 61.725 ;
        RECT 109.940 61.555 110.110 61.725 ;
        RECT 110.300 61.555 110.470 61.725 ;
        RECT 110.660 61.555 110.830 61.725 ;
        RECT 111.020 61.555 111.190 61.725 ;
        RECT 111.380 61.555 111.550 61.725 ;
        RECT 112.220 61.555 112.390 61.725 ;
        RECT 112.580 61.555 112.750 61.725 ;
        RECT 112.940 61.555 113.110 61.725 ;
        RECT 113.300 61.555 113.470 61.725 ;
        RECT 113.660 61.555 113.830 61.725 ;
        RECT 114.500 61.555 114.670 61.725 ;
        RECT 114.860 61.555 115.030 61.725 ;
        RECT 115.220 61.555 115.390 61.725 ;
        RECT 115.580 61.555 115.750 61.725 ;
        RECT 115.940 61.555 116.110 61.725 ;
        RECT 116.780 61.555 116.950 61.725 ;
        RECT 117.140 61.555 117.310 61.725 ;
        RECT 117.500 61.555 117.670 61.725 ;
        RECT 117.860 61.555 118.030 61.725 ;
        RECT 118.220 61.555 118.390 61.725 ;
        RECT 119.060 61.555 119.230 61.725 ;
        RECT 119.420 61.555 119.590 61.725 ;
        RECT 119.780 61.555 119.950 61.725 ;
        RECT 120.140 61.555 120.310 61.725 ;
        RECT 120.500 61.555 120.670 61.725 ;
        RECT 121.340 61.555 121.510 61.725 ;
        RECT 121.700 61.555 121.870 61.725 ;
        RECT 122.060 61.555 122.230 61.725 ;
        RECT 122.420 61.555 122.590 61.725 ;
        RECT 122.780 61.555 122.950 61.725 ;
        RECT 123.620 61.555 123.790 61.725 ;
        RECT 123.980 61.555 124.150 61.725 ;
        RECT 124.340 61.555 124.510 61.725 ;
        RECT 124.700 61.555 124.870 61.725 ;
        RECT 125.060 61.555 125.230 61.725 ;
        RECT 125.900 61.555 126.070 61.725 ;
        RECT 126.260 61.555 126.430 61.725 ;
        RECT 126.620 61.555 126.790 61.725 ;
        RECT 126.980 61.555 127.150 61.725 ;
        RECT 127.340 61.555 127.510 61.725 ;
        RECT 128.180 61.555 128.350 61.725 ;
        RECT 128.540 61.555 128.710 61.725 ;
        RECT 128.900 61.555 129.070 61.725 ;
        RECT 129.260 61.555 129.430 61.725 ;
        RECT 129.620 61.555 129.790 61.725 ;
        RECT 130.460 61.555 130.630 61.725 ;
        RECT 130.820 61.555 130.990 61.725 ;
        RECT 131.180 61.555 131.350 61.725 ;
        RECT 131.540 61.555 131.710 61.725 ;
        RECT 131.900 61.555 132.070 61.725 ;
        RECT 132.740 61.555 132.910 61.725 ;
        RECT 133.100 61.555 133.270 61.725 ;
        RECT 133.460 61.555 133.630 61.725 ;
        RECT 133.820 61.555 133.990 61.725 ;
        RECT 134.180 61.555 134.350 61.725 ;
        RECT 135.020 61.555 135.190 61.725 ;
        RECT 135.380 61.555 135.550 61.725 ;
        RECT 135.740 61.555 135.910 61.725 ;
        RECT 136.100 61.555 136.270 61.725 ;
        RECT 136.460 61.555 136.630 61.725 ;
        RECT 137.300 61.555 137.470 61.725 ;
        RECT 137.660 61.555 137.830 61.725 ;
        RECT 138.020 61.555 138.190 61.725 ;
        RECT 138.380 61.555 138.550 61.725 ;
        RECT 138.740 61.555 138.910 61.725 ;
        RECT 139.580 61.555 139.750 61.725 ;
        RECT 139.940 61.555 140.110 61.725 ;
        RECT 140.300 61.555 140.470 61.725 ;
        RECT 140.660 61.555 140.830 61.725 ;
        RECT 141.020 61.555 141.190 61.725 ;
        RECT 141.860 61.555 142.030 61.725 ;
        RECT 142.220 61.555 142.390 61.725 ;
        RECT 142.580 61.555 142.750 61.725 ;
        RECT 142.940 61.555 143.110 61.725 ;
        RECT 143.300 61.555 143.470 61.725 ;
        RECT 144.390 61.495 144.560 61.665 ;
        RECT 42.730 61.185 42.900 61.355 ;
        RECT 33.580 60.690 33.750 60.860 ;
        RECT 33.580 60.330 33.750 60.500 ;
        RECT 34.500 60.445 34.670 60.615 ;
        RECT 34.860 60.445 35.030 60.615 ;
        RECT 35.360 60.445 35.530 60.615 ;
        RECT 35.720 60.445 35.890 60.615 ;
        RECT 36.220 60.445 36.390 60.615 ;
        RECT 36.580 60.445 36.750 60.615 ;
        RECT 37.080 60.445 37.250 60.615 ;
        RECT 37.440 60.445 37.610 60.615 ;
        RECT 38.360 60.690 38.530 60.860 ;
        RECT 38.360 60.330 38.530 60.500 ;
        RECT 33.580 59.970 33.750 60.140 ;
        RECT 33.580 59.610 33.750 59.780 ;
        RECT 33.580 59.250 33.750 59.420 ;
        RECT 34.250 59.790 34.420 59.960 ;
        RECT 34.250 59.430 34.420 59.600 ;
        RECT 34.680 59.790 34.850 59.960 ;
        RECT 34.680 59.430 34.850 59.600 ;
        RECT 35.110 59.790 35.280 59.960 ;
        RECT 35.110 59.430 35.280 59.600 ;
        RECT 35.540 59.790 35.710 59.960 ;
        RECT 35.540 59.430 35.710 59.600 ;
        RECT 35.970 59.790 36.140 59.960 ;
        RECT 35.970 59.430 36.140 59.600 ;
        RECT 36.400 59.790 36.570 59.960 ;
        RECT 36.400 59.430 36.570 59.600 ;
        RECT 36.830 59.790 37.000 59.960 ;
        RECT 36.830 59.430 37.000 59.600 ;
        RECT 37.260 59.790 37.430 59.960 ;
        RECT 37.260 59.430 37.430 59.600 ;
        RECT 37.690 59.790 37.860 59.960 ;
        RECT 37.690 59.430 37.860 59.600 ;
        RECT 38.360 59.970 38.530 60.140 ;
        RECT 38.360 59.610 38.530 59.780 ;
        RECT 42.730 60.825 42.900 60.995 ;
        RECT 42.730 60.465 42.900 60.635 ;
        RECT 43.400 61.050 43.570 61.220 ;
        RECT 43.400 60.690 43.570 60.860 ;
        RECT 45.680 61.050 45.850 61.220 ;
        RECT 45.680 60.690 45.850 60.860 ;
        RECT 47.960 61.050 48.130 61.220 ;
        RECT 47.960 60.690 48.130 60.860 ;
        RECT 50.240 61.050 50.410 61.220 ;
        RECT 50.240 60.690 50.410 60.860 ;
        RECT 52.520 61.050 52.690 61.220 ;
        RECT 52.520 60.690 52.690 60.860 ;
        RECT 54.800 61.050 54.970 61.220 ;
        RECT 54.800 60.690 54.970 60.860 ;
        RECT 57.080 61.050 57.250 61.220 ;
        RECT 57.080 60.690 57.250 60.860 ;
        RECT 59.360 61.050 59.530 61.220 ;
        RECT 59.360 60.690 59.530 60.860 ;
        RECT 61.640 61.050 61.810 61.220 ;
        RECT 61.640 60.690 61.810 60.860 ;
        RECT 63.920 61.050 64.090 61.220 ;
        RECT 63.920 60.690 64.090 60.860 ;
        RECT 66.200 61.050 66.370 61.220 ;
        RECT 66.200 60.690 66.370 60.860 ;
        RECT 68.480 61.050 68.650 61.220 ;
        RECT 68.480 60.690 68.650 60.860 ;
        RECT 70.760 61.050 70.930 61.220 ;
        RECT 70.760 60.690 70.930 60.860 ;
        RECT 73.040 61.050 73.210 61.220 ;
        RECT 73.040 60.690 73.210 60.860 ;
        RECT 75.320 61.050 75.490 61.220 ;
        RECT 75.320 60.690 75.490 60.860 ;
        RECT 77.600 61.050 77.770 61.220 ;
        RECT 77.600 60.690 77.770 60.860 ;
        RECT 79.880 61.050 80.050 61.220 ;
        RECT 79.880 60.690 80.050 60.860 ;
        RECT 82.160 61.050 82.330 61.220 ;
        RECT 82.160 60.690 82.330 60.860 ;
        RECT 84.440 61.050 84.610 61.220 ;
        RECT 84.440 60.690 84.610 60.860 ;
        RECT 86.720 61.050 86.890 61.220 ;
        RECT 86.720 60.690 86.890 60.860 ;
        RECT 89.000 61.050 89.170 61.220 ;
        RECT 89.000 60.690 89.170 60.860 ;
        RECT 91.280 61.050 91.450 61.220 ;
        RECT 91.280 60.690 91.450 60.860 ;
        RECT 93.560 61.050 93.730 61.220 ;
        RECT 93.560 60.690 93.730 60.860 ;
        RECT 95.840 61.050 96.010 61.220 ;
        RECT 95.840 60.690 96.010 60.860 ;
        RECT 98.120 61.050 98.290 61.220 ;
        RECT 98.120 60.690 98.290 60.860 ;
        RECT 100.400 61.050 100.570 61.220 ;
        RECT 100.400 60.690 100.570 60.860 ;
        RECT 102.680 61.050 102.850 61.220 ;
        RECT 102.680 60.690 102.850 60.860 ;
        RECT 104.960 61.050 105.130 61.220 ;
        RECT 104.960 60.690 105.130 60.860 ;
        RECT 107.240 61.050 107.410 61.220 ;
        RECT 107.240 60.690 107.410 60.860 ;
        RECT 109.520 61.050 109.690 61.220 ;
        RECT 109.520 60.690 109.690 60.860 ;
        RECT 111.800 61.050 111.970 61.220 ;
        RECT 111.800 60.690 111.970 60.860 ;
        RECT 114.080 61.050 114.250 61.220 ;
        RECT 114.080 60.690 114.250 60.860 ;
        RECT 116.360 61.050 116.530 61.220 ;
        RECT 116.360 60.690 116.530 60.860 ;
        RECT 118.640 61.050 118.810 61.220 ;
        RECT 118.640 60.690 118.810 60.860 ;
        RECT 120.920 61.050 121.090 61.220 ;
        RECT 120.920 60.690 121.090 60.860 ;
        RECT 123.200 61.050 123.370 61.220 ;
        RECT 123.200 60.690 123.370 60.860 ;
        RECT 125.480 61.050 125.650 61.220 ;
        RECT 125.480 60.690 125.650 60.860 ;
        RECT 127.760 61.050 127.930 61.220 ;
        RECT 127.760 60.690 127.930 60.860 ;
        RECT 130.040 61.050 130.210 61.220 ;
        RECT 130.040 60.690 130.210 60.860 ;
        RECT 132.320 61.050 132.490 61.220 ;
        RECT 132.320 60.690 132.490 60.860 ;
        RECT 134.600 61.050 134.770 61.220 ;
        RECT 134.600 60.690 134.770 60.860 ;
        RECT 136.880 61.050 137.050 61.220 ;
        RECT 136.880 60.690 137.050 60.860 ;
        RECT 139.160 61.050 139.330 61.220 ;
        RECT 139.160 60.690 139.330 60.860 ;
        RECT 141.440 61.050 141.610 61.220 ;
        RECT 141.440 60.690 141.610 60.860 ;
        RECT 143.720 61.050 143.890 61.220 ;
        RECT 143.720 60.690 143.890 60.860 ;
        RECT 144.390 61.135 144.560 61.305 ;
        RECT 144.390 60.775 144.560 60.945 ;
        RECT 42.730 60.105 42.900 60.275 ;
        RECT 144.390 60.415 144.560 60.585 ;
        RECT 144.390 60.055 144.560 60.225 ;
        RECT 42.790 59.635 42.960 59.805 ;
        RECT 43.150 59.635 43.320 59.805 ;
        RECT 43.510 59.635 43.680 59.805 ;
        RECT 43.870 59.635 44.040 59.805 ;
        RECT 44.230 59.635 44.400 59.805 ;
        RECT 44.590 59.635 44.760 59.805 ;
        RECT 44.950 59.635 45.120 59.805 ;
        RECT 45.310 59.635 45.480 59.805 ;
        RECT 45.670 59.635 45.840 59.805 ;
        RECT 46.030 59.635 46.200 59.805 ;
        RECT 46.390 59.635 46.560 59.805 ;
        RECT 46.750 59.635 46.920 59.805 ;
        RECT 47.110 59.635 47.280 59.805 ;
        RECT 47.470 59.635 47.640 59.805 ;
        RECT 47.830 59.635 48.000 59.805 ;
        RECT 48.190 59.635 48.360 59.805 ;
        RECT 48.550 59.635 48.720 59.805 ;
        RECT 48.910 59.635 49.080 59.805 ;
        RECT 49.270 59.635 49.440 59.805 ;
        RECT 49.630 59.635 49.800 59.805 ;
        RECT 49.990 59.635 50.160 59.805 ;
        RECT 50.350 59.635 50.520 59.805 ;
        RECT 50.710 59.635 50.880 59.805 ;
        RECT 51.070 59.635 51.240 59.805 ;
        RECT 51.430 59.635 51.600 59.805 ;
        RECT 51.790 59.635 51.960 59.805 ;
        RECT 52.150 59.635 52.320 59.805 ;
        RECT 52.510 59.635 52.680 59.805 ;
        RECT 52.870 59.635 53.040 59.805 ;
        RECT 53.230 59.635 53.400 59.805 ;
        RECT 53.590 59.635 53.760 59.805 ;
        RECT 53.950 59.635 54.120 59.805 ;
        RECT 54.310 59.635 54.480 59.805 ;
        RECT 54.670 59.635 54.840 59.805 ;
        RECT 55.030 59.635 55.200 59.805 ;
        RECT 55.390 59.635 55.560 59.805 ;
        RECT 55.750 59.635 55.920 59.805 ;
        RECT 56.110 59.635 56.280 59.805 ;
        RECT 56.470 59.635 56.640 59.805 ;
        RECT 56.830 59.635 57.000 59.805 ;
        RECT 57.190 59.635 57.360 59.805 ;
        RECT 57.550 59.635 57.720 59.805 ;
        RECT 57.910 59.635 58.080 59.805 ;
        RECT 58.270 59.635 58.440 59.805 ;
        RECT 58.630 59.635 58.800 59.805 ;
        RECT 58.990 59.635 59.160 59.805 ;
        RECT 59.350 59.635 59.520 59.805 ;
        RECT 59.710 59.635 59.880 59.805 ;
        RECT 60.070 59.635 60.240 59.805 ;
        RECT 60.430 59.635 60.600 59.805 ;
        RECT 60.790 59.635 60.960 59.805 ;
        RECT 61.150 59.635 61.320 59.805 ;
        RECT 61.510 59.635 61.680 59.805 ;
        RECT 61.870 59.635 62.040 59.805 ;
        RECT 62.230 59.635 62.400 59.805 ;
        RECT 62.590 59.635 62.760 59.805 ;
        RECT 62.950 59.635 63.120 59.805 ;
        RECT 63.310 59.635 63.480 59.805 ;
        RECT 63.670 59.635 63.840 59.805 ;
        RECT 64.030 59.635 64.200 59.805 ;
        RECT 64.390 59.635 64.560 59.805 ;
        RECT 64.750 59.635 64.920 59.805 ;
        RECT 65.110 59.635 65.280 59.805 ;
        RECT 65.470 59.635 65.640 59.805 ;
        RECT 65.830 59.635 66.000 59.805 ;
        RECT 66.190 59.635 66.360 59.805 ;
        RECT 66.550 59.635 66.720 59.805 ;
        RECT 66.910 59.635 67.080 59.805 ;
        RECT 67.270 59.635 67.440 59.805 ;
        RECT 67.630 59.635 67.800 59.805 ;
        RECT 67.990 59.635 68.160 59.805 ;
        RECT 68.350 59.635 68.520 59.805 ;
        RECT 68.710 59.635 68.880 59.805 ;
        RECT 69.070 59.635 69.240 59.805 ;
        RECT 69.430 59.635 69.600 59.805 ;
        RECT 69.790 59.635 69.960 59.805 ;
        RECT 70.150 59.635 70.320 59.805 ;
        RECT 70.510 59.635 70.680 59.805 ;
        RECT 70.870 59.635 71.040 59.805 ;
        RECT 71.230 59.635 71.400 59.805 ;
        RECT 71.590 59.635 71.760 59.805 ;
        RECT 71.950 59.635 72.120 59.805 ;
        RECT 72.310 59.635 72.480 59.805 ;
        RECT 72.670 59.635 72.840 59.805 ;
        RECT 73.030 59.635 73.200 59.805 ;
        RECT 73.390 59.635 73.560 59.805 ;
        RECT 73.750 59.635 73.920 59.805 ;
        RECT 74.110 59.635 74.280 59.805 ;
        RECT 74.470 59.635 74.640 59.805 ;
        RECT 74.830 59.635 75.000 59.805 ;
        RECT 75.190 59.635 75.360 59.805 ;
        RECT 75.550 59.635 75.720 59.805 ;
        RECT 75.910 59.635 76.080 59.805 ;
        RECT 76.270 59.635 76.440 59.805 ;
        RECT 76.630 59.635 76.800 59.805 ;
        RECT 76.990 59.635 77.160 59.805 ;
        RECT 77.350 59.635 77.520 59.805 ;
        RECT 77.710 59.635 77.880 59.805 ;
        RECT 78.070 59.635 78.240 59.805 ;
        RECT 78.430 59.635 78.600 59.805 ;
        RECT 78.790 59.635 78.960 59.805 ;
        RECT 79.150 59.635 79.320 59.805 ;
        RECT 79.510 59.635 79.680 59.805 ;
        RECT 79.870 59.635 80.040 59.805 ;
        RECT 80.230 59.635 80.400 59.805 ;
        RECT 80.590 59.635 80.760 59.805 ;
        RECT 80.950 59.635 81.120 59.805 ;
        RECT 81.310 59.635 81.480 59.805 ;
        RECT 81.670 59.635 81.840 59.805 ;
        RECT 82.030 59.635 82.200 59.805 ;
        RECT 82.390 59.635 82.560 59.805 ;
        RECT 82.750 59.635 82.920 59.805 ;
        RECT 83.110 59.635 83.280 59.805 ;
        RECT 83.470 59.635 83.640 59.805 ;
        RECT 83.830 59.635 84.000 59.805 ;
        RECT 84.190 59.635 84.360 59.805 ;
        RECT 84.550 59.635 84.720 59.805 ;
        RECT 84.910 59.635 85.080 59.805 ;
        RECT 85.270 59.635 85.440 59.805 ;
        RECT 85.630 59.635 85.800 59.805 ;
        RECT 85.990 59.635 86.160 59.805 ;
        RECT 86.350 59.635 86.520 59.805 ;
        RECT 86.710 59.635 86.880 59.805 ;
        RECT 87.070 59.635 87.240 59.805 ;
        RECT 87.430 59.635 87.600 59.805 ;
        RECT 87.790 59.635 87.960 59.805 ;
        RECT 88.150 59.635 88.320 59.805 ;
        RECT 88.510 59.635 88.680 59.805 ;
        RECT 88.870 59.635 89.040 59.805 ;
        RECT 89.230 59.635 89.400 59.805 ;
        RECT 89.590 59.635 89.760 59.805 ;
        RECT 89.950 59.635 90.120 59.805 ;
        RECT 90.310 59.635 90.480 59.805 ;
        RECT 90.670 59.635 90.840 59.805 ;
        RECT 91.030 59.635 91.200 59.805 ;
        RECT 91.390 59.635 91.560 59.805 ;
        RECT 91.750 59.635 91.920 59.805 ;
        RECT 92.110 59.635 92.280 59.805 ;
        RECT 92.470 59.635 92.640 59.805 ;
        RECT 92.830 59.635 93.000 59.805 ;
        RECT 93.190 59.635 93.360 59.805 ;
        RECT 93.740 59.635 93.910 59.805 ;
        RECT 94.100 59.635 94.270 59.805 ;
        RECT 94.460 59.635 94.630 59.805 ;
        RECT 94.820 59.635 94.990 59.805 ;
        RECT 95.180 59.635 95.350 59.805 ;
        RECT 95.540 59.635 95.710 59.805 ;
        RECT 95.900 59.635 96.070 59.805 ;
        RECT 96.260 59.635 96.430 59.805 ;
        RECT 96.620 59.635 96.790 59.805 ;
        RECT 96.980 59.635 97.150 59.805 ;
        RECT 97.340 59.635 97.510 59.805 ;
        RECT 97.700 59.635 97.870 59.805 ;
        RECT 98.060 59.635 98.230 59.805 ;
        RECT 98.420 59.635 98.590 59.805 ;
        RECT 98.780 59.635 98.950 59.805 ;
        RECT 99.140 59.635 99.310 59.805 ;
        RECT 99.500 59.635 99.670 59.805 ;
        RECT 99.860 59.635 100.030 59.805 ;
        RECT 100.220 59.635 100.390 59.805 ;
        RECT 100.580 59.635 100.750 59.805 ;
        RECT 100.940 59.635 101.110 59.805 ;
        RECT 101.300 59.635 101.470 59.805 ;
        RECT 101.660 59.635 101.830 59.805 ;
        RECT 102.020 59.635 102.190 59.805 ;
        RECT 102.380 59.635 102.550 59.805 ;
        RECT 102.740 59.635 102.910 59.805 ;
        RECT 103.100 59.635 103.270 59.805 ;
        RECT 103.460 59.635 103.630 59.805 ;
        RECT 103.820 59.635 103.990 59.805 ;
        RECT 104.180 59.635 104.350 59.805 ;
        RECT 104.540 59.635 104.710 59.805 ;
        RECT 104.900 59.635 105.070 59.805 ;
        RECT 105.260 59.635 105.430 59.805 ;
        RECT 105.620 59.635 105.790 59.805 ;
        RECT 105.980 59.635 106.150 59.805 ;
        RECT 106.340 59.635 106.510 59.805 ;
        RECT 106.700 59.635 106.870 59.805 ;
        RECT 107.060 59.635 107.230 59.805 ;
        RECT 107.420 59.635 107.590 59.805 ;
        RECT 107.780 59.635 107.950 59.805 ;
        RECT 108.140 59.635 108.310 59.805 ;
        RECT 108.500 59.635 108.670 59.805 ;
        RECT 108.860 59.635 109.030 59.805 ;
        RECT 109.220 59.635 109.390 59.805 ;
        RECT 109.580 59.635 109.750 59.805 ;
        RECT 109.940 59.635 110.110 59.805 ;
        RECT 110.300 59.635 110.470 59.805 ;
        RECT 110.660 59.635 110.830 59.805 ;
        RECT 111.020 59.635 111.190 59.805 ;
        RECT 111.380 59.635 111.550 59.805 ;
        RECT 111.740 59.635 111.910 59.805 ;
        RECT 112.100 59.635 112.270 59.805 ;
        RECT 112.460 59.635 112.630 59.805 ;
        RECT 112.820 59.635 112.990 59.805 ;
        RECT 113.180 59.635 113.350 59.805 ;
        RECT 113.540 59.635 113.710 59.805 ;
        RECT 113.900 59.635 114.070 59.805 ;
        RECT 114.260 59.635 114.430 59.805 ;
        RECT 114.620 59.635 114.790 59.805 ;
        RECT 114.980 59.635 115.150 59.805 ;
        RECT 115.340 59.635 115.510 59.805 ;
        RECT 115.700 59.635 115.870 59.805 ;
        RECT 116.060 59.635 116.230 59.805 ;
        RECT 116.420 59.635 116.590 59.805 ;
        RECT 116.780 59.635 116.950 59.805 ;
        RECT 117.140 59.635 117.310 59.805 ;
        RECT 117.500 59.635 117.670 59.805 ;
        RECT 117.860 59.635 118.030 59.805 ;
        RECT 118.220 59.635 118.390 59.805 ;
        RECT 118.580 59.635 118.750 59.805 ;
        RECT 118.940 59.635 119.110 59.805 ;
        RECT 119.300 59.635 119.470 59.805 ;
        RECT 119.660 59.635 119.830 59.805 ;
        RECT 120.020 59.635 120.190 59.805 ;
        RECT 120.380 59.635 120.550 59.805 ;
        RECT 120.740 59.635 120.910 59.805 ;
        RECT 121.100 59.635 121.270 59.805 ;
        RECT 121.460 59.635 121.630 59.805 ;
        RECT 121.820 59.635 121.990 59.805 ;
        RECT 122.180 59.635 122.350 59.805 ;
        RECT 122.540 59.635 122.710 59.805 ;
        RECT 122.900 59.635 123.070 59.805 ;
        RECT 123.260 59.635 123.430 59.805 ;
        RECT 123.620 59.635 123.790 59.805 ;
        RECT 123.980 59.635 124.150 59.805 ;
        RECT 124.340 59.635 124.510 59.805 ;
        RECT 124.700 59.635 124.870 59.805 ;
        RECT 125.060 59.635 125.230 59.805 ;
        RECT 125.420 59.635 125.590 59.805 ;
        RECT 125.780 59.635 125.950 59.805 ;
        RECT 126.140 59.635 126.310 59.805 ;
        RECT 126.500 59.635 126.670 59.805 ;
        RECT 126.860 59.635 127.030 59.805 ;
        RECT 127.220 59.635 127.390 59.805 ;
        RECT 127.580 59.635 127.750 59.805 ;
        RECT 127.940 59.635 128.110 59.805 ;
        RECT 128.300 59.635 128.470 59.805 ;
        RECT 128.660 59.635 128.830 59.805 ;
        RECT 129.020 59.635 129.190 59.805 ;
        RECT 129.380 59.635 129.550 59.805 ;
        RECT 129.740 59.635 129.910 59.805 ;
        RECT 130.100 59.635 130.270 59.805 ;
        RECT 130.460 59.635 130.630 59.805 ;
        RECT 130.820 59.635 130.990 59.805 ;
        RECT 131.180 59.635 131.350 59.805 ;
        RECT 131.540 59.635 131.710 59.805 ;
        RECT 131.900 59.635 132.070 59.805 ;
        RECT 132.260 59.635 132.430 59.805 ;
        RECT 132.620 59.635 132.790 59.805 ;
        RECT 132.980 59.635 133.150 59.805 ;
        RECT 133.340 59.635 133.510 59.805 ;
        RECT 133.700 59.635 133.870 59.805 ;
        RECT 134.060 59.635 134.230 59.805 ;
        RECT 134.420 59.635 134.590 59.805 ;
        RECT 134.780 59.635 134.950 59.805 ;
        RECT 135.140 59.635 135.310 59.805 ;
        RECT 135.500 59.635 135.670 59.805 ;
        RECT 135.860 59.635 136.030 59.805 ;
        RECT 136.220 59.635 136.390 59.805 ;
        RECT 136.580 59.635 136.750 59.805 ;
        RECT 136.940 59.635 137.110 59.805 ;
        RECT 137.300 59.635 137.470 59.805 ;
        RECT 137.660 59.635 137.830 59.805 ;
        RECT 138.020 59.635 138.190 59.805 ;
        RECT 138.380 59.635 138.550 59.805 ;
        RECT 138.740 59.635 138.910 59.805 ;
        RECT 139.100 59.635 139.270 59.805 ;
        RECT 139.460 59.635 139.630 59.805 ;
        RECT 139.820 59.635 139.990 59.805 ;
        RECT 140.180 59.635 140.350 59.805 ;
        RECT 140.540 59.635 140.710 59.805 ;
        RECT 140.900 59.635 141.070 59.805 ;
        RECT 141.260 59.635 141.430 59.805 ;
        RECT 141.620 59.635 141.790 59.805 ;
        RECT 141.980 59.635 142.150 59.805 ;
        RECT 142.340 59.635 142.510 59.805 ;
        RECT 142.700 59.635 142.870 59.805 ;
        RECT 143.060 59.635 143.230 59.805 ;
        RECT 143.420 59.635 143.590 59.805 ;
        RECT 143.780 59.635 143.950 59.805 ;
        RECT 144.390 59.695 144.560 59.865 ;
        RECT 38.360 59.250 38.530 59.420 ;
        RECT 33.580 58.890 33.750 59.060 ;
        RECT 38.360 58.890 38.530 59.060 ;
        RECT 33.930 58.590 34.100 58.760 ;
        RECT 34.290 58.590 34.460 58.760 ;
        RECT 34.650 58.590 34.820 58.760 ;
        RECT 35.010 58.590 35.180 58.760 ;
        RECT 35.370 58.590 35.540 58.760 ;
        RECT 35.730 58.590 35.900 58.760 ;
        RECT 36.090 58.590 36.260 58.760 ;
        RECT 36.450 58.590 36.620 58.760 ;
        RECT 36.810 58.590 36.980 58.760 ;
        RECT 37.170 58.590 37.340 58.760 ;
        RECT 37.530 58.590 37.700 58.760 ;
        RECT 37.890 58.590 38.060 58.760 ;
        RECT 56.330 53.440 56.500 53.610 ;
        RECT 56.690 53.440 56.860 53.610 ;
        RECT 57.050 53.440 57.220 53.610 ;
        RECT 57.410 53.440 57.580 53.610 ;
        RECT 57.770 53.440 57.940 53.610 ;
        RECT 58.130 53.440 58.300 53.610 ;
        RECT 58.490 53.440 58.660 53.610 ;
        RECT 58.850 53.440 59.020 53.610 ;
        RECT 59.210 53.440 59.380 53.610 ;
        RECT 59.570 53.440 59.740 53.610 ;
        RECT 59.930 53.440 60.100 53.610 ;
        RECT 60.290 53.440 60.460 53.610 ;
        RECT 60.650 53.440 60.820 53.610 ;
        RECT 61.010 53.440 61.180 53.610 ;
        RECT 61.370 53.440 61.540 53.610 ;
        RECT 61.730 53.440 61.900 53.610 ;
        RECT 62.090 53.440 62.260 53.610 ;
        RECT 62.450 53.440 62.620 53.610 ;
        RECT 62.810 53.440 62.980 53.610 ;
        RECT 63.170 53.440 63.340 53.610 ;
        RECT 63.530 53.440 63.700 53.610 ;
        RECT 63.890 53.440 64.060 53.610 ;
        RECT 64.250 53.440 64.420 53.610 ;
        RECT 64.610 53.440 64.780 53.610 ;
        RECT 64.970 53.440 65.140 53.610 ;
        RECT 65.330 53.440 65.500 53.610 ;
        RECT 65.690 53.440 65.860 53.610 ;
        RECT 66.050 53.440 66.220 53.610 ;
        RECT 66.410 53.440 66.580 53.610 ;
        RECT 66.770 53.440 66.940 53.610 ;
        RECT 67.130 53.440 67.300 53.610 ;
        RECT 67.490 53.440 67.660 53.610 ;
        RECT 67.850 53.440 68.020 53.610 ;
        RECT 68.210 53.440 68.380 53.610 ;
        RECT 68.570 53.440 68.740 53.610 ;
        RECT 68.930 53.440 69.100 53.610 ;
        RECT 69.290 53.440 69.460 53.610 ;
        RECT 69.650 53.440 69.820 53.610 ;
        RECT 70.010 53.440 70.180 53.610 ;
        RECT 70.370 53.440 70.540 53.610 ;
        RECT 70.730 53.440 70.900 53.610 ;
        RECT 71.090 53.440 71.260 53.610 ;
        RECT 71.450 53.440 71.620 53.610 ;
        RECT 71.810 53.440 71.980 53.610 ;
        RECT 72.170 53.440 72.340 53.610 ;
        RECT 72.530 53.440 72.700 53.610 ;
        RECT 72.890 53.440 73.060 53.610 ;
        RECT 73.250 53.440 73.420 53.610 ;
        RECT 73.610 53.440 73.780 53.610 ;
        RECT 73.970 53.440 74.140 53.610 ;
        RECT 74.330 53.440 74.500 53.610 ;
        RECT 74.690 53.440 74.860 53.610 ;
        RECT 75.050 53.440 75.220 53.610 ;
        RECT 75.410 53.440 75.580 53.610 ;
        RECT 75.770 53.440 75.940 53.610 ;
        RECT 76.130 53.440 76.300 53.610 ;
        RECT 76.490 53.440 76.660 53.610 ;
        RECT 76.850 53.440 77.020 53.610 ;
        RECT 77.210 53.440 77.380 53.610 ;
        RECT 77.570 53.440 77.740 53.610 ;
        RECT 77.930 53.440 78.100 53.610 ;
        RECT 78.290 53.440 78.460 53.610 ;
        RECT 78.650 53.440 78.820 53.610 ;
        RECT 79.010 53.440 79.180 53.610 ;
        RECT 79.370 53.440 79.540 53.610 ;
        RECT 79.730 53.440 79.900 53.610 ;
        RECT 80.090 53.440 80.260 53.610 ;
        RECT 80.450 53.440 80.620 53.610 ;
        RECT 80.810 53.440 80.980 53.610 ;
        RECT 81.170 53.440 81.340 53.610 ;
        RECT 81.530 53.440 81.700 53.610 ;
        RECT 81.890 53.440 82.060 53.610 ;
        RECT 82.250 53.440 82.420 53.610 ;
        RECT 82.610 53.440 82.780 53.610 ;
        RECT 82.970 53.440 83.140 53.610 ;
        RECT 83.330 53.440 83.500 53.610 ;
        RECT 83.690 53.440 83.860 53.610 ;
        RECT 84.050 53.440 84.220 53.610 ;
        RECT 84.410 53.440 84.580 53.610 ;
        RECT 84.770 53.440 84.940 53.610 ;
        RECT 85.130 53.440 85.300 53.610 ;
        RECT 85.490 53.440 85.660 53.610 ;
        RECT 85.850 53.440 86.020 53.610 ;
        RECT 86.210 53.440 86.380 53.610 ;
        RECT 86.570 53.440 86.740 53.610 ;
        RECT 86.930 53.440 87.100 53.610 ;
        RECT 87.290 53.440 87.460 53.610 ;
        RECT 87.650 53.440 87.820 53.610 ;
        RECT 88.010 53.440 88.180 53.610 ;
        RECT 88.370 53.440 88.540 53.610 ;
        RECT 88.730 53.440 88.900 53.610 ;
        RECT 89.090 53.440 89.260 53.610 ;
        RECT 89.450 53.440 89.620 53.610 ;
        RECT 89.810 53.440 89.980 53.610 ;
        RECT 90.170 53.440 90.340 53.610 ;
        RECT 90.530 53.440 90.700 53.610 ;
        RECT 90.890 53.440 91.060 53.610 ;
        RECT 91.250 53.440 91.420 53.610 ;
        RECT 91.610 53.440 91.780 53.610 ;
        RECT 91.970 53.440 92.140 53.610 ;
        RECT 92.330 53.440 92.500 53.610 ;
        RECT 92.690 53.440 92.860 53.610 ;
        RECT 93.050 53.440 93.220 53.610 ;
        RECT 93.410 53.440 93.580 53.610 ;
        RECT 93.770 53.440 93.940 53.610 ;
        RECT 94.130 53.440 94.300 53.610 ;
        RECT 94.490 53.440 94.660 53.610 ;
        RECT 94.850 53.440 95.020 53.610 ;
        RECT 55.980 53.140 56.150 53.310 ;
        RECT 95.480 53.140 95.650 53.310 ;
        RECT 55.980 52.780 56.150 52.950 ;
        RECT 77.710 52.890 77.880 53.060 ;
        RECT 78.070 52.890 78.240 53.060 ;
        RECT 78.430 52.890 78.600 53.060 ;
        RECT 78.790 52.890 78.960 53.060 ;
        RECT 79.150 52.890 79.320 53.060 ;
        RECT 79.990 52.890 80.160 53.060 ;
        RECT 80.350 52.890 80.520 53.060 ;
        RECT 80.710 52.890 80.880 53.060 ;
        RECT 81.070 52.890 81.240 53.060 ;
        RECT 81.430 52.890 81.600 53.060 ;
        RECT 95.480 52.780 95.650 52.950 ;
        RECT 55.980 52.420 56.150 52.590 ;
        RECT 55.980 52.060 56.150 52.230 ;
        RECT 55.980 51.700 56.150 51.870 ;
        RECT 65.890 52.235 66.060 52.405 ;
        RECT 65.890 51.875 66.060 52.045 ;
        RECT 68.170 52.235 68.340 52.405 ;
        RECT 68.170 51.875 68.340 52.045 ;
        RECT 70.450 52.235 70.620 52.405 ;
        RECT 70.450 51.875 70.620 52.045 ;
        RECT 72.730 52.235 72.900 52.405 ;
        RECT 72.730 51.875 72.900 52.045 ;
        RECT 75.010 52.235 75.180 52.405 ;
        RECT 75.010 51.875 75.180 52.045 ;
        RECT 77.290 52.235 77.460 52.405 ;
        RECT 77.290 51.875 77.460 52.045 ;
        RECT 79.570 52.235 79.740 52.405 ;
        RECT 79.570 51.875 79.740 52.045 ;
        RECT 81.850 52.235 82.020 52.405 ;
        RECT 81.850 51.875 82.020 52.045 ;
        RECT 84.130 52.235 84.300 52.405 ;
        RECT 84.130 51.875 84.300 52.045 ;
        RECT 86.410 52.235 86.580 52.405 ;
        RECT 86.410 51.875 86.580 52.045 ;
        RECT 88.690 52.235 88.860 52.405 ;
        RECT 88.690 51.875 88.860 52.045 ;
        RECT 90.970 52.235 91.140 52.405 ;
        RECT 90.970 51.875 91.140 52.045 ;
        RECT 93.250 52.235 93.420 52.405 ;
        RECT 93.250 51.875 93.420 52.045 ;
        RECT 95.480 52.420 95.650 52.590 ;
        RECT 95.480 52.060 95.650 52.230 ;
        RECT 95.480 51.700 95.650 51.870 ;
        RECT 55.980 51.340 56.150 51.510 ;
        RECT 55.980 50.980 56.150 51.150 ;
        RECT 66.310 51.220 66.480 51.390 ;
        RECT 66.670 51.220 66.840 51.390 ;
        RECT 67.030 51.220 67.200 51.390 ;
        RECT 67.390 51.220 67.560 51.390 ;
        RECT 67.750 51.220 67.920 51.390 ;
        RECT 68.590 51.220 68.760 51.390 ;
        RECT 68.950 51.220 69.120 51.390 ;
        RECT 69.310 51.220 69.480 51.390 ;
        RECT 69.670 51.220 69.840 51.390 ;
        RECT 70.030 51.220 70.200 51.390 ;
        RECT 70.870 51.220 71.040 51.390 ;
        RECT 71.230 51.220 71.400 51.390 ;
        RECT 71.590 51.220 71.760 51.390 ;
        RECT 71.950 51.220 72.120 51.390 ;
        RECT 72.310 51.220 72.480 51.390 ;
        RECT 73.150 51.220 73.320 51.390 ;
        RECT 73.510 51.220 73.680 51.390 ;
        RECT 73.870 51.220 74.040 51.390 ;
        RECT 74.230 51.220 74.400 51.390 ;
        RECT 74.590 51.220 74.760 51.390 ;
        RECT 75.430 51.220 75.600 51.390 ;
        RECT 75.790 51.220 75.960 51.390 ;
        RECT 76.150 51.220 76.320 51.390 ;
        RECT 76.510 51.220 76.680 51.390 ;
        RECT 76.870 51.220 77.040 51.390 ;
        RECT 82.270 51.220 82.440 51.390 ;
        RECT 82.630 51.220 82.800 51.390 ;
        RECT 82.990 51.220 83.160 51.390 ;
        RECT 83.350 51.220 83.520 51.390 ;
        RECT 83.710 51.220 83.880 51.390 ;
        RECT 84.550 51.220 84.720 51.390 ;
        RECT 84.910 51.220 85.080 51.390 ;
        RECT 85.270 51.220 85.440 51.390 ;
        RECT 85.630 51.220 85.800 51.390 ;
        RECT 85.990 51.220 86.160 51.390 ;
        RECT 86.830 51.220 87.000 51.390 ;
        RECT 87.190 51.220 87.360 51.390 ;
        RECT 87.550 51.220 87.720 51.390 ;
        RECT 87.910 51.220 88.080 51.390 ;
        RECT 88.270 51.220 88.440 51.390 ;
        RECT 89.110 51.220 89.280 51.390 ;
        RECT 89.470 51.220 89.640 51.390 ;
        RECT 89.830 51.220 90.000 51.390 ;
        RECT 90.190 51.220 90.360 51.390 ;
        RECT 90.550 51.220 90.720 51.390 ;
        RECT 91.390 51.220 91.560 51.390 ;
        RECT 91.750 51.220 91.920 51.390 ;
        RECT 92.110 51.220 92.280 51.390 ;
        RECT 92.470 51.220 92.640 51.390 ;
        RECT 92.830 51.220 93.000 51.390 ;
        RECT 95.480 51.340 95.650 51.510 ;
        RECT 55.980 50.620 56.150 50.790 ;
        RECT 55.980 50.260 56.150 50.430 ;
        RECT 55.980 49.900 56.150 50.070 ;
        RECT 55.980 49.540 56.150 49.710 ;
        RECT 95.480 50.980 95.650 51.150 ;
        RECT 95.480 50.620 95.650 50.790 ;
        RECT 95.480 50.260 95.650 50.430 ;
        RECT 95.480 49.900 95.650 50.070 ;
        RECT 55.980 49.180 56.150 49.350 ;
        RECT 57.070 49.300 57.240 49.470 ;
        RECT 57.430 49.300 57.600 49.470 ;
        RECT 57.790 49.300 57.960 49.470 ;
        RECT 63.190 49.300 63.360 49.470 ;
        RECT 63.550 49.300 63.720 49.470 ;
        RECT 63.910 49.300 64.080 49.470 ;
        RECT 64.750 49.300 64.920 49.470 ;
        RECT 65.110 49.300 65.280 49.470 ;
        RECT 65.470 49.300 65.640 49.470 ;
        RECT 66.310 49.300 66.480 49.470 ;
        RECT 66.670 49.300 66.840 49.470 ;
        RECT 67.030 49.300 67.200 49.470 ;
        RECT 67.390 49.300 67.560 49.470 ;
        RECT 67.750 49.300 67.920 49.470 ;
        RECT 68.590 49.300 68.760 49.470 ;
        RECT 68.950 49.300 69.120 49.470 ;
        RECT 69.310 49.300 69.480 49.470 ;
        RECT 69.670 49.300 69.840 49.470 ;
        RECT 70.030 49.300 70.200 49.470 ;
        RECT 70.870 49.300 71.040 49.470 ;
        RECT 71.230 49.300 71.400 49.470 ;
        RECT 71.590 49.300 71.760 49.470 ;
        RECT 71.950 49.300 72.120 49.470 ;
        RECT 72.310 49.300 72.480 49.470 ;
        RECT 73.150 49.300 73.320 49.470 ;
        RECT 73.510 49.300 73.680 49.470 ;
        RECT 73.870 49.300 74.040 49.470 ;
        RECT 74.230 49.300 74.400 49.470 ;
        RECT 74.590 49.300 74.760 49.470 ;
        RECT 75.430 49.300 75.600 49.470 ;
        RECT 75.790 49.300 75.960 49.470 ;
        RECT 76.150 49.300 76.320 49.470 ;
        RECT 76.510 49.300 76.680 49.470 ;
        RECT 76.870 49.300 77.040 49.470 ;
        RECT 77.710 49.300 77.880 49.470 ;
        RECT 78.070 49.300 78.240 49.470 ;
        RECT 78.430 49.300 78.600 49.470 ;
        RECT 78.790 49.300 78.960 49.470 ;
        RECT 79.150 49.300 79.320 49.470 ;
        RECT 79.990 49.300 80.160 49.470 ;
        RECT 80.350 49.300 80.520 49.470 ;
        RECT 80.710 49.300 80.880 49.470 ;
        RECT 81.070 49.300 81.240 49.470 ;
        RECT 81.430 49.300 81.600 49.470 ;
        RECT 82.270 49.300 82.440 49.470 ;
        RECT 82.630 49.300 82.800 49.470 ;
        RECT 82.990 49.300 83.160 49.470 ;
        RECT 83.350 49.300 83.520 49.470 ;
        RECT 83.710 49.300 83.880 49.470 ;
        RECT 84.550 49.300 84.720 49.470 ;
        RECT 84.910 49.300 85.080 49.470 ;
        RECT 85.270 49.300 85.440 49.470 ;
        RECT 85.630 49.300 85.800 49.470 ;
        RECT 85.990 49.300 86.160 49.470 ;
        RECT 86.830 49.300 87.000 49.470 ;
        RECT 87.190 49.300 87.360 49.470 ;
        RECT 87.550 49.300 87.720 49.470 ;
        RECT 87.910 49.300 88.080 49.470 ;
        RECT 88.270 49.300 88.440 49.470 ;
        RECT 89.110 49.300 89.280 49.470 ;
        RECT 89.470 49.300 89.640 49.470 ;
        RECT 89.830 49.300 90.000 49.470 ;
        RECT 90.190 49.300 90.360 49.470 ;
        RECT 90.550 49.300 90.720 49.470 ;
        RECT 91.390 49.300 91.560 49.470 ;
        RECT 91.750 49.300 91.920 49.470 ;
        RECT 92.110 49.300 92.280 49.470 ;
        RECT 92.470 49.300 92.640 49.470 ;
        RECT 92.830 49.300 93.000 49.470 ;
        RECT 93.670 49.300 93.840 49.470 ;
        RECT 94.030 49.300 94.200 49.470 ;
        RECT 94.390 49.300 94.560 49.470 ;
        RECT 95.480 49.540 95.650 49.710 ;
        RECT 95.480 49.180 95.650 49.350 ;
        RECT 55.980 48.820 56.150 48.990 ;
        RECT 55.980 48.460 56.150 48.630 ;
        RECT 55.980 48.100 56.150 48.270 ;
        RECT 56.650 48.645 56.820 48.815 ;
        RECT 56.650 48.285 56.820 48.455 ;
        RECT 57.430 48.645 57.600 48.815 ;
        RECT 57.430 48.285 57.600 48.455 ;
        RECT 58.210 48.645 58.380 48.815 ;
        RECT 58.210 48.285 58.380 48.455 ;
        RECT 60.490 48.645 60.660 48.815 ;
        RECT 60.490 48.285 60.660 48.455 ;
        RECT 62.770 48.645 62.940 48.815 ;
        RECT 62.770 48.285 62.940 48.455 ;
        RECT 63.550 48.645 63.720 48.815 ;
        RECT 63.550 48.285 63.720 48.455 ;
        RECT 64.330 48.645 64.500 48.815 ;
        RECT 64.330 48.285 64.500 48.455 ;
        RECT 65.110 48.645 65.280 48.815 ;
        RECT 65.110 48.285 65.280 48.455 ;
        RECT 65.890 48.645 66.060 48.815 ;
        RECT 65.890 48.285 66.060 48.455 ;
        RECT 68.170 48.645 68.340 48.815 ;
        RECT 68.170 48.285 68.340 48.455 ;
        RECT 70.450 48.645 70.620 48.815 ;
        RECT 70.450 48.285 70.620 48.455 ;
        RECT 72.730 48.645 72.900 48.815 ;
        RECT 72.730 48.285 72.900 48.455 ;
        RECT 75.010 48.645 75.180 48.815 ;
        RECT 75.010 48.285 75.180 48.455 ;
        RECT 77.290 48.645 77.460 48.815 ;
        RECT 77.290 48.285 77.460 48.455 ;
        RECT 79.570 48.645 79.740 48.815 ;
        RECT 79.570 48.285 79.740 48.455 ;
        RECT 81.850 48.645 82.020 48.815 ;
        RECT 81.850 48.285 82.020 48.455 ;
        RECT 84.130 48.645 84.300 48.815 ;
        RECT 84.130 48.285 84.300 48.455 ;
        RECT 86.410 48.645 86.580 48.815 ;
        RECT 86.410 48.285 86.580 48.455 ;
        RECT 88.690 48.645 88.860 48.815 ;
        RECT 88.690 48.285 88.860 48.455 ;
        RECT 90.970 48.645 91.140 48.815 ;
        RECT 90.970 48.285 91.140 48.455 ;
        RECT 93.250 48.645 93.420 48.815 ;
        RECT 93.250 48.285 93.420 48.455 ;
        RECT 94.030 48.645 94.200 48.815 ;
        RECT 94.030 48.285 94.200 48.455 ;
        RECT 94.810 48.645 94.980 48.815 ;
        RECT 94.810 48.285 94.980 48.455 ;
        RECT 95.480 48.820 95.650 48.990 ;
        RECT 95.480 48.460 95.650 48.630 ;
        RECT 95.480 48.100 95.650 48.270 ;
        RECT 55.980 47.740 56.150 47.910 ;
        RECT 58.630 47.630 58.800 47.800 ;
        RECT 58.990 47.630 59.160 47.800 ;
        RECT 59.350 47.630 59.520 47.800 ;
        RECT 59.710 47.630 59.880 47.800 ;
        RECT 60.070 47.630 60.240 47.800 ;
        RECT 60.910 47.630 61.080 47.800 ;
        RECT 61.270 47.630 61.440 47.800 ;
        RECT 61.630 47.630 61.800 47.800 ;
        RECT 61.990 47.630 62.160 47.800 ;
        RECT 62.350 47.630 62.520 47.800 ;
        RECT 66.310 47.630 66.480 47.800 ;
        RECT 66.670 47.630 66.840 47.800 ;
        RECT 67.030 47.630 67.200 47.800 ;
        RECT 67.390 47.630 67.560 47.800 ;
        RECT 67.750 47.630 67.920 47.800 ;
        RECT 68.590 47.630 68.760 47.800 ;
        RECT 68.950 47.630 69.120 47.800 ;
        RECT 69.310 47.630 69.480 47.800 ;
        RECT 69.670 47.630 69.840 47.800 ;
        RECT 70.030 47.630 70.200 47.800 ;
        RECT 70.870 47.630 71.040 47.800 ;
        RECT 71.230 47.630 71.400 47.800 ;
        RECT 71.590 47.630 71.760 47.800 ;
        RECT 71.950 47.630 72.120 47.800 ;
        RECT 72.310 47.630 72.480 47.800 ;
        RECT 73.150 47.630 73.320 47.800 ;
        RECT 73.510 47.630 73.680 47.800 ;
        RECT 73.870 47.630 74.040 47.800 ;
        RECT 74.230 47.630 74.400 47.800 ;
        RECT 74.590 47.630 74.760 47.800 ;
        RECT 75.430 47.630 75.600 47.800 ;
        RECT 75.790 47.630 75.960 47.800 ;
        RECT 76.150 47.630 76.320 47.800 ;
        RECT 76.510 47.630 76.680 47.800 ;
        RECT 76.870 47.630 77.040 47.800 ;
        RECT 77.710 47.630 77.880 47.800 ;
        RECT 78.070 47.630 78.240 47.800 ;
        RECT 78.430 47.630 78.600 47.800 ;
        RECT 78.790 47.630 78.960 47.800 ;
        RECT 79.150 47.630 79.320 47.800 ;
        RECT 79.990 47.630 80.160 47.800 ;
        RECT 80.350 47.630 80.520 47.800 ;
        RECT 80.710 47.630 80.880 47.800 ;
        RECT 81.070 47.630 81.240 47.800 ;
        RECT 81.430 47.630 81.600 47.800 ;
        RECT 82.270 47.630 82.440 47.800 ;
        RECT 82.630 47.630 82.800 47.800 ;
        RECT 82.990 47.630 83.160 47.800 ;
        RECT 83.350 47.630 83.520 47.800 ;
        RECT 83.710 47.630 83.880 47.800 ;
        RECT 84.550 47.630 84.720 47.800 ;
        RECT 84.910 47.630 85.080 47.800 ;
        RECT 85.270 47.630 85.440 47.800 ;
        RECT 85.630 47.630 85.800 47.800 ;
        RECT 85.990 47.630 86.160 47.800 ;
        RECT 86.830 47.630 87.000 47.800 ;
        RECT 87.190 47.630 87.360 47.800 ;
        RECT 87.550 47.630 87.720 47.800 ;
        RECT 87.910 47.630 88.080 47.800 ;
        RECT 88.270 47.630 88.440 47.800 ;
        RECT 89.110 47.630 89.280 47.800 ;
        RECT 89.470 47.630 89.640 47.800 ;
        RECT 89.830 47.630 90.000 47.800 ;
        RECT 90.190 47.630 90.360 47.800 ;
        RECT 90.550 47.630 90.720 47.800 ;
        RECT 91.390 47.630 91.560 47.800 ;
        RECT 91.750 47.630 91.920 47.800 ;
        RECT 92.110 47.630 92.280 47.800 ;
        RECT 92.470 47.630 92.640 47.800 ;
        RECT 92.830 47.630 93.000 47.800 ;
        RECT 95.480 47.740 95.650 47.910 ;
        RECT 55.980 47.380 56.150 47.550 ;
        RECT 95.480 47.380 95.650 47.550 ;
        RECT 56.330 47.080 56.500 47.250 ;
        RECT 56.690 47.080 56.860 47.250 ;
        RECT 57.050 47.080 57.220 47.250 ;
        RECT 57.410 47.080 57.580 47.250 ;
        RECT 57.770 47.080 57.940 47.250 ;
        RECT 58.130 47.080 58.300 47.250 ;
        RECT 58.490 47.080 58.660 47.250 ;
        RECT 58.850 47.080 59.020 47.250 ;
        RECT 59.210 47.080 59.380 47.250 ;
        RECT 59.570 47.080 59.740 47.250 ;
        RECT 59.930 47.080 60.100 47.250 ;
        RECT 60.290 47.080 60.460 47.250 ;
        RECT 60.650 47.080 60.820 47.250 ;
        RECT 61.010 47.080 61.180 47.250 ;
        RECT 61.370 47.080 61.540 47.250 ;
        RECT 61.730 47.080 61.900 47.250 ;
        RECT 62.090 47.080 62.260 47.250 ;
        RECT 62.450 47.080 62.620 47.250 ;
        RECT 62.810 47.080 62.980 47.250 ;
        RECT 63.170 47.080 63.340 47.250 ;
        RECT 63.530 47.080 63.700 47.250 ;
        RECT 63.890 47.080 64.060 47.250 ;
        RECT 64.250 47.080 64.420 47.250 ;
        RECT 64.610 47.080 64.780 47.250 ;
        RECT 64.970 47.080 65.140 47.250 ;
        RECT 65.330 47.080 65.500 47.250 ;
        RECT 65.690 47.080 65.860 47.250 ;
        RECT 66.050 47.080 66.220 47.250 ;
        RECT 66.410 47.080 66.580 47.250 ;
        RECT 66.770 47.080 66.940 47.250 ;
        RECT 67.130 47.080 67.300 47.250 ;
        RECT 67.490 47.080 67.660 47.250 ;
        RECT 67.850 47.080 68.020 47.250 ;
        RECT 68.210 47.080 68.380 47.250 ;
        RECT 68.570 47.080 68.740 47.250 ;
        RECT 68.930 47.080 69.100 47.250 ;
        RECT 69.290 47.080 69.460 47.250 ;
        RECT 69.650 47.080 69.820 47.250 ;
        RECT 70.010 47.080 70.180 47.250 ;
        RECT 70.370 47.080 70.540 47.250 ;
        RECT 70.730 47.080 70.900 47.250 ;
        RECT 71.090 47.080 71.260 47.250 ;
        RECT 71.450 47.080 71.620 47.250 ;
        RECT 71.810 47.080 71.980 47.250 ;
        RECT 72.170 47.080 72.340 47.250 ;
        RECT 72.530 47.080 72.700 47.250 ;
        RECT 72.890 47.080 73.060 47.250 ;
        RECT 73.250 47.080 73.420 47.250 ;
        RECT 73.610 47.080 73.780 47.250 ;
        RECT 73.970 47.080 74.140 47.250 ;
        RECT 74.330 47.080 74.500 47.250 ;
        RECT 74.690 47.080 74.860 47.250 ;
        RECT 75.050 47.080 75.220 47.250 ;
        RECT 75.410 47.080 75.580 47.250 ;
        RECT 75.770 47.080 75.940 47.250 ;
        RECT 76.130 47.080 76.300 47.250 ;
        RECT 76.490 47.080 76.660 47.250 ;
        RECT 76.850 47.080 77.020 47.250 ;
        RECT 77.210 47.080 77.380 47.250 ;
        RECT 77.570 47.080 77.740 47.250 ;
        RECT 77.930 47.080 78.100 47.250 ;
        RECT 78.290 47.080 78.460 47.250 ;
        RECT 78.650 47.080 78.820 47.250 ;
        RECT 79.010 47.080 79.180 47.250 ;
        RECT 79.370 47.080 79.540 47.250 ;
        RECT 79.730 47.080 79.900 47.250 ;
        RECT 80.090 47.080 80.260 47.250 ;
        RECT 80.450 47.080 80.620 47.250 ;
        RECT 80.810 47.080 80.980 47.250 ;
        RECT 81.170 47.080 81.340 47.250 ;
        RECT 81.530 47.080 81.700 47.250 ;
        RECT 81.890 47.080 82.060 47.250 ;
        RECT 82.250 47.080 82.420 47.250 ;
        RECT 82.610 47.080 82.780 47.250 ;
        RECT 82.970 47.080 83.140 47.250 ;
        RECT 83.330 47.080 83.500 47.250 ;
        RECT 83.690 47.080 83.860 47.250 ;
        RECT 84.050 47.080 84.220 47.250 ;
        RECT 84.410 47.080 84.580 47.250 ;
        RECT 84.770 47.080 84.940 47.250 ;
        RECT 85.130 47.080 85.300 47.250 ;
        RECT 85.490 47.080 85.660 47.250 ;
        RECT 85.850 47.080 86.020 47.250 ;
        RECT 86.210 47.080 86.380 47.250 ;
        RECT 86.570 47.080 86.740 47.250 ;
        RECT 86.930 47.080 87.100 47.250 ;
        RECT 87.290 47.080 87.460 47.250 ;
        RECT 87.650 47.080 87.820 47.250 ;
        RECT 88.010 47.080 88.180 47.250 ;
        RECT 88.370 47.080 88.540 47.250 ;
        RECT 88.730 47.080 88.900 47.250 ;
        RECT 89.090 47.080 89.260 47.250 ;
        RECT 89.450 47.080 89.620 47.250 ;
        RECT 89.810 47.080 89.980 47.250 ;
        RECT 90.170 47.080 90.340 47.250 ;
        RECT 90.530 47.080 90.700 47.250 ;
        RECT 90.890 47.080 91.060 47.250 ;
        RECT 91.250 47.080 91.420 47.250 ;
        RECT 91.610 47.080 91.780 47.250 ;
        RECT 91.970 47.080 92.140 47.250 ;
        RECT 92.330 47.080 92.500 47.250 ;
        RECT 92.690 47.080 92.860 47.250 ;
        RECT 93.050 47.080 93.220 47.250 ;
        RECT 93.410 47.080 93.580 47.250 ;
        RECT 93.770 47.080 93.940 47.250 ;
        RECT 94.130 47.080 94.300 47.250 ;
        RECT 94.490 47.080 94.660 47.250 ;
        RECT 94.850 47.080 95.020 47.250 ;
        RECT 94.490 45.935 94.660 46.105 ;
        RECT 94.850 45.935 95.020 46.105 ;
        RECT 95.210 45.935 95.380 46.105 ;
        RECT 95.570 45.935 95.740 46.105 ;
        RECT 95.930 45.935 96.100 46.105 ;
        RECT 96.290 45.935 96.460 46.105 ;
        RECT 96.650 45.935 96.820 46.105 ;
        RECT 97.010 45.935 97.180 46.105 ;
        RECT 97.370 45.935 97.540 46.105 ;
        RECT 97.730 45.935 97.900 46.105 ;
        RECT 98.090 45.935 98.260 46.105 ;
        RECT 98.450 45.935 98.620 46.105 ;
        RECT 98.810 45.935 98.980 46.105 ;
        RECT 99.170 45.935 99.340 46.105 ;
        RECT 99.530 45.935 99.700 46.105 ;
        RECT 99.890 45.935 100.060 46.105 ;
        RECT 100.250 45.935 100.420 46.105 ;
        RECT 100.610 45.935 100.780 46.105 ;
        RECT 100.970 45.935 101.140 46.105 ;
        RECT 101.330 45.935 101.500 46.105 ;
        RECT 101.690 45.935 101.860 46.105 ;
        RECT 102.050 45.935 102.220 46.105 ;
        RECT 102.410 45.935 102.580 46.105 ;
        RECT 102.770 45.935 102.940 46.105 ;
        RECT 103.130 45.935 103.300 46.105 ;
        RECT 103.490 45.935 103.660 46.105 ;
        RECT 103.850 45.935 104.020 46.105 ;
        RECT 104.210 45.935 104.380 46.105 ;
        RECT 104.570 45.935 104.740 46.105 ;
        RECT 104.930 45.935 105.100 46.105 ;
        RECT 105.290 45.935 105.460 46.105 ;
        RECT 105.650 45.935 105.820 46.105 ;
        RECT 106.010 45.935 106.180 46.105 ;
        RECT 106.370 45.935 106.540 46.105 ;
        RECT 106.730 45.935 106.900 46.105 ;
        RECT 107.090 45.935 107.260 46.105 ;
        RECT 107.450 45.935 107.620 46.105 ;
        RECT 107.810 45.935 107.980 46.105 ;
        RECT 108.170 45.935 108.340 46.105 ;
        RECT 108.530 45.935 108.700 46.105 ;
        RECT 108.890 45.935 109.060 46.105 ;
        RECT 109.250 45.935 109.420 46.105 ;
        RECT 109.610 45.935 109.780 46.105 ;
        RECT 109.970 45.935 110.140 46.105 ;
        RECT 110.330 45.935 110.500 46.105 ;
        RECT 110.690 45.935 110.860 46.105 ;
        RECT 111.050 45.935 111.220 46.105 ;
        RECT 111.410 45.935 111.580 46.105 ;
        RECT 111.770 45.935 111.940 46.105 ;
        RECT 112.130 45.935 112.300 46.105 ;
        RECT 112.490 45.935 112.660 46.105 ;
        RECT 112.850 45.935 113.020 46.105 ;
        RECT 113.210 45.935 113.380 46.105 ;
        RECT 113.570 45.935 113.740 46.105 ;
        RECT 113.930 45.935 114.100 46.105 ;
        RECT 114.290 45.935 114.460 46.105 ;
        RECT 114.650 45.935 114.820 46.105 ;
        RECT 115.010 45.935 115.180 46.105 ;
        RECT 115.370 45.935 115.540 46.105 ;
        RECT 115.730 45.935 115.900 46.105 ;
        RECT 116.090 45.935 116.260 46.105 ;
        RECT 116.450 45.935 116.620 46.105 ;
        RECT 116.810 45.935 116.980 46.105 ;
        RECT 117.170 45.935 117.340 46.105 ;
        RECT 117.530 45.935 117.700 46.105 ;
        RECT 117.890 45.935 118.060 46.105 ;
        RECT 94.140 45.635 94.310 45.805 ;
        RECT 118.280 45.635 118.450 45.805 ;
        RECT 56.330 45.185 56.500 45.355 ;
        RECT 56.690 45.185 56.860 45.355 ;
        RECT 57.050 45.185 57.220 45.355 ;
        RECT 57.410 45.185 57.580 45.355 ;
        RECT 57.770 45.185 57.940 45.355 ;
        RECT 58.130 45.185 58.300 45.355 ;
        RECT 58.490 45.185 58.660 45.355 ;
        RECT 58.850 45.185 59.020 45.355 ;
        RECT 59.210 45.185 59.380 45.355 ;
        RECT 59.570 45.185 59.740 45.355 ;
        RECT 59.930 45.185 60.100 45.355 ;
        RECT 60.290 45.185 60.460 45.355 ;
        RECT 60.650 45.185 60.820 45.355 ;
        RECT 61.010 45.185 61.180 45.355 ;
        RECT 61.370 45.185 61.540 45.355 ;
        RECT 61.730 45.185 61.900 45.355 ;
        RECT 62.090 45.185 62.260 45.355 ;
        RECT 62.450 45.185 62.620 45.355 ;
        RECT 62.810 45.185 62.980 45.355 ;
        RECT 63.170 45.185 63.340 45.355 ;
        RECT 63.530 45.185 63.700 45.355 ;
        RECT 63.890 45.185 64.060 45.355 ;
        RECT 64.250 45.185 64.420 45.355 ;
        RECT 64.610 45.185 64.780 45.355 ;
        RECT 55.980 44.655 56.150 44.825 ;
        RECT 58.630 44.635 58.800 44.805 ;
        RECT 58.990 44.635 59.160 44.805 ;
        RECT 59.350 44.635 59.520 44.805 ;
        RECT 59.710 44.635 59.880 44.805 ;
        RECT 60.070 44.635 60.240 44.805 ;
        RECT 60.910 44.635 61.080 44.805 ;
        RECT 61.270 44.635 61.440 44.805 ;
        RECT 61.630 44.635 61.800 44.805 ;
        RECT 61.990 44.635 62.160 44.805 ;
        RECT 62.350 44.635 62.520 44.805 ;
        RECT 65.000 44.655 65.170 44.825 ;
        RECT 55.980 44.295 56.150 44.465 ;
        RECT 55.980 43.935 56.150 44.105 ;
        RECT 56.650 44.050 56.820 44.220 ;
        RECT 57.430 44.050 57.600 44.220 ;
        RECT 58.210 44.050 58.380 44.220 ;
        RECT 60.490 44.050 60.660 44.220 ;
        RECT 62.770 44.050 62.940 44.220 ;
        RECT 63.550 44.050 63.720 44.220 ;
        RECT 64.330 44.050 64.500 44.220 ;
        RECT 65.000 44.295 65.170 44.465 ;
        RECT 65.000 43.935 65.170 44.105 ;
        RECT 55.980 43.575 56.150 43.745 ;
        RECT 57.070 43.465 57.240 43.635 ;
        RECT 57.430 43.465 57.600 43.635 ;
        RECT 57.790 43.465 57.960 43.635 ;
        RECT 63.190 43.465 63.360 43.635 ;
        RECT 63.550 43.465 63.720 43.635 ;
        RECT 63.910 43.465 64.080 43.635 ;
        RECT 65.000 43.575 65.170 43.745 ;
        RECT 55.980 43.215 56.150 43.385 ;
        RECT 65.000 43.215 65.170 43.385 ;
        RECT 56.330 42.915 56.500 43.085 ;
        RECT 56.690 42.915 56.860 43.085 ;
        RECT 57.050 42.915 57.220 43.085 ;
        RECT 57.410 42.915 57.580 43.085 ;
        RECT 57.770 42.915 57.940 43.085 ;
        RECT 58.130 42.915 58.300 43.085 ;
        RECT 58.490 42.915 58.660 43.085 ;
        RECT 58.850 42.915 59.020 43.085 ;
        RECT 59.210 42.915 59.380 43.085 ;
        RECT 59.570 42.915 59.740 43.085 ;
        RECT 59.930 42.915 60.100 43.085 ;
        RECT 60.290 42.915 60.460 43.085 ;
        RECT 60.650 42.915 60.820 43.085 ;
        RECT 61.010 42.915 61.180 43.085 ;
        RECT 61.370 42.915 61.540 43.085 ;
        RECT 61.730 42.915 61.900 43.085 ;
        RECT 62.090 42.915 62.260 43.085 ;
        RECT 62.450 42.915 62.620 43.085 ;
        RECT 62.810 42.915 62.980 43.085 ;
        RECT 63.170 42.915 63.340 43.085 ;
        RECT 63.530 42.915 63.700 43.085 ;
        RECT 63.890 42.915 64.060 43.085 ;
        RECT 64.250 42.915 64.420 43.085 ;
        RECT 64.610 42.915 64.780 43.085 ;
        RECT 69.540 45.185 69.710 45.355 ;
        RECT 69.900 45.185 70.070 45.355 ;
        RECT 70.260 45.185 70.430 45.355 ;
        RECT 70.620 45.185 70.790 45.355 ;
        RECT 70.980 45.185 71.150 45.355 ;
        RECT 71.340 45.185 71.510 45.355 ;
        RECT 71.700 45.185 71.870 45.355 ;
        RECT 72.060 45.185 72.230 45.355 ;
        RECT 72.420 45.185 72.590 45.355 ;
        RECT 72.780 45.185 72.950 45.355 ;
        RECT 73.140 45.185 73.310 45.355 ;
        RECT 73.500 45.185 73.670 45.355 ;
        RECT 73.860 45.185 74.030 45.355 ;
        RECT 74.220 45.185 74.390 45.355 ;
        RECT 74.580 45.185 74.750 45.355 ;
        RECT 74.940 45.185 75.110 45.355 ;
        RECT 75.300 45.185 75.470 45.355 ;
        RECT 75.660 45.185 75.830 45.355 ;
        RECT 76.020 45.185 76.190 45.355 ;
        RECT 76.380 45.185 76.550 45.355 ;
        RECT 76.740 45.185 76.910 45.355 ;
        RECT 77.100 45.185 77.270 45.355 ;
        RECT 77.460 45.185 77.630 45.355 ;
        RECT 77.820 45.185 77.990 45.355 ;
        RECT 78.180 45.185 78.350 45.355 ;
        RECT 78.540 45.185 78.710 45.355 ;
        RECT 78.900 45.185 79.070 45.355 ;
        RECT 79.260 45.185 79.430 45.355 ;
        RECT 79.620 45.185 79.790 45.355 ;
        RECT 79.980 45.185 80.150 45.355 ;
        RECT 80.340 45.185 80.510 45.355 ;
        RECT 80.700 45.185 80.870 45.355 ;
        RECT 81.060 45.185 81.230 45.355 ;
        RECT 81.420 45.185 81.590 45.355 ;
        RECT 81.780 45.185 81.950 45.355 ;
        RECT 82.140 45.185 82.310 45.355 ;
        RECT 82.500 45.185 82.670 45.355 ;
        RECT 82.860 45.185 83.030 45.355 ;
        RECT 83.220 45.185 83.390 45.355 ;
        RECT 83.580 45.185 83.750 45.355 ;
        RECT 83.940 45.185 84.110 45.355 ;
        RECT 84.300 45.185 84.470 45.355 ;
        RECT 84.660 45.185 84.830 45.355 ;
        RECT 85.020 45.185 85.190 45.355 ;
        RECT 85.380 45.185 85.550 45.355 ;
        RECT 85.740 45.185 85.910 45.355 ;
        RECT 86.100 45.185 86.270 45.355 ;
        RECT 86.460 45.185 86.630 45.355 ;
        RECT 86.820 45.185 86.990 45.355 ;
        RECT 87.180 45.185 87.350 45.355 ;
        RECT 87.540 45.185 87.710 45.355 ;
        RECT 87.900 45.185 88.070 45.355 ;
        RECT 88.260 45.185 88.430 45.355 ;
        RECT 88.620 45.185 88.790 45.355 ;
        RECT 88.980 45.185 89.150 45.355 ;
        RECT 89.340 45.185 89.510 45.355 ;
        RECT 69.190 44.655 69.360 44.825 ;
        RECT 70.245 44.635 70.415 44.805 ;
        RECT 70.605 44.635 70.775 44.805 ;
        RECT 70.965 44.635 71.135 44.805 ;
        RECT 71.325 44.635 71.495 44.805 ;
        RECT 71.685 44.635 71.855 44.805 ;
        RECT 72.045 44.635 72.215 44.805 ;
        RECT 72.840 44.635 73.010 44.805 ;
        RECT 73.200 44.635 73.370 44.805 ;
        RECT 73.560 44.635 73.730 44.805 ;
        RECT 73.920 44.635 74.090 44.805 ;
        RECT 74.280 44.635 74.450 44.805 ;
        RECT 75.120 44.635 75.290 44.805 ;
        RECT 75.480 44.635 75.650 44.805 ;
        RECT 75.840 44.635 76.010 44.805 ;
        RECT 76.200 44.635 76.370 44.805 ;
        RECT 76.560 44.635 76.730 44.805 ;
        RECT 77.365 44.635 77.535 44.805 ;
        RECT 77.725 44.635 77.895 44.805 ;
        RECT 78.085 44.635 78.255 44.805 ;
        RECT 78.445 44.635 78.615 44.805 ;
        RECT 78.805 44.635 78.975 44.805 ;
        RECT 79.165 44.635 79.335 44.805 ;
        RECT 79.925 44.635 80.095 44.805 ;
        RECT 80.285 44.635 80.455 44.805 ;
        RECT 80.645 44.635 80.815 44.805 ;
        RECT 81.005 44.635 81.175 44.805 ;
        RECT 81.365 44.635 81.535 44.805 ;
        RECT 81.725 44.635 81.895 44.805 ;
        RECT 82.520 44.635 82.690 44.805 ;
        RECT 82.880 44.635 83.050 44.805 ;
        RECT 83.240 44.635 83.410 44.805 ;
        RECT 83.600 44.635 83.770 44.805 ;
        RECT 83.960 44.635 84.130 44.805 ;
        RECT 84.800 44.635 84.970 44.805 ;
        RECT 85.160 44.635 85.330 44.805 ;
        RECT 85.520 44.635 85.690 44.805 ;
        RECT 85.880 44.635 86.050 44.805 ;
        RECT 86.240 44.635 86.410 44.805 ;
        RECT 87.045 44.635 87.215 44.805 ;
        RECT 87.405 44.635 87.575 44.805 ;
        RECT 87.765 44.635 87.935 44.805 ;
        RECT 88.125 44.635 88.295 44.805 ;
        RECT 88.485 44.635 88.655 44.805 ;
        RECT 88.845 44.635 89.015 44.805 ;
        RECT 89.890 44.655 90.060 44.825 ;
        RECT 69.190 44.295 69.360 44.465 ;
        RECT 69.190 43.935 69.360 44.105 ;
        RECT 69.860 44.050 70.030 44.220 ;
        RECT 71.140 44.050 71.310 44.220 ;
        RECT 72.420 44.050 72.590 44.220 ;
        RECT 74.700 44.050 74.870 44.220 ;
        RECT 76.980 44.050 77.150 44.220 ;
        RECT 78.260 44.050 78.430 44.220 ;
        RECT 79.540 44.050 79.710 44.220 ;
        RECT 80.820 44.050 80.990 44.220 ;
        RECT 82.100 44.050 82.270 44.220 ;
        RECT 84.380 44.050 84.550 44.220 ;
        RECT 86.660 44.050 86.830 44.220 ;
        RECT 87.940 44.050 88.110 44.220 ;
        RECT 89.220 44.050 89.390 44.220 ;
        RECT 89.890 44.295 90.060 44.465 ;
        RECT 89.890 43.935 90.060 44.105 ;
        RECT 69.190 43.575 69.360 43.745 ;
        RECT 70.245 43.465 70.415 43.635 ;
        RECT 70.605 43.465 70.775 43.635 ;
        RECT 70.965 43.465 71.135 43.635 ;
        RECT 71.325 43.465 71.495 43.635 ;
        RECT 71.685 43.465 71.855 43.635 ;
        RECT 72.045 43.465 72.215 43.635 ;
        RECT 72.840 43.465 73.010 43.635 ;
        RECT 73.200 43.465 73.370 43.635 ;
        RECT 73.560 43.465 73.730 43.635 ;
        RECT 73.920 43.465 74.090 43.635 ;
        RECT 74.280 43.465 74.450 43.635 ;
        RECT 75.120 43.465 75.290 43.635 ;
        RECT 75.480 43.465 75.650 43.635 ;
        RECT 75.840 43.465 76.010 43.635 ;
        RECT 76.200 43.465 76.370 43.635 ;
        RECT 76.560 43.465 76.730 43.635 ;
        RECT 77.365 43.465 77.535 43.635 ;
        RECT 77.725 43.465 77.895 43.635 ;
        RECT 78.085 43.465 78.255 43.635 ;
        RECT 78.445 43.465 78.615 43.635 ;
        RECT 78.805 43.465 78.975 43.635 ;
        RECT 79.165 43.465 79.335 43.635 ;
        RECT 79.925 43.465 80.095 43.635 ;
        RECT 80.285 43.465 80.455 43.635 ;
        RECT 80.645 43.465 80.815 43.635 ;
        RECT 81.005 43.465 81.175 43.635 ;
        RECT 81.365 43.465 81.535 43.635 ;
        RECT 81.725 43.465 81.895 43.635 ;
        RECT 87.045 43.465 87.215 43.635 ;
        RECT 87.405 43.465 87.575 43.635 ;
        RECT 87.765 43.465 87.935 43.635 ;
        RECT 88.125 43.465 88.295 43.635 ;
        RECT 88.485 43.465 88.655 43.635 ;
        RECT 88.845 43.465 89.015 43.635 ;
        RECT 89.890 43.575 90.060 43.745 ;
        RECT 69.190 43.215 69.360 43.385 ;
        RECT 89.890 43.215 90.060 43.385 ;
        RECT 69.540 42.915 69.710 43.085 ;
        RECT 69.900 42.915 70.070 43.085 ;
        RECT 70.260 42.915 70.430 43.085 ;
        RECT 70.620 42.915 70.790 43.085 ;
        RECT 70.980 42.915 71.150 43.085 ;
        RECT 71.340 42.915 71.510 43.085 ;
        RECT 71.700 42.915 71.870 43.085 ;
        RECT 72.060 42.915 72.230 43.085 ;
        RECT 72.420 42.915 72.590 43.085 ;
        RECT 72.780 42.915 72.950 43.085 ;
        RECT 73.140 42.915 73.310 43.085 ;
        RECT 73.500 42.915 73.670 43.085 ;
        RECT 73.860 42.915 74.030 43.085 ;
        RECT 74.220 42.915 74.390 43.085 ;
        RECT 74.580 42.915 74.750 43.085 ;
        RECT 74.940 42.915 75.110 43.085 ;
        RECT 75.300 42.915 75.470 43.085 ;
        RECT 75.660 42.915 75.830 43.085 ;
        RECT 76.020 42.915 76.190 43.085 ;
        RECT 76.380 42.915 76.550 43.085 ;
        RECT 76.740 42.915 76.910 43.085 ;
        RECT 77.100 42.915 77.270 43.085 ;
        RECT 77.460 42.915 77.630 43.085 ;
        RECT 77.820 42.915 77.990 43.085 ;
        RECT 78.180 42.915 78.350 43.085 ;
        RECT 78.540 42.915 78.710 43.085 ;
        RECT 78.900 42.915 79.070 43.085 ;
        RECT 79.260 42.915 79.430 43.085 ;
        RECT 79.620 42.915 79.790 43.085 ;
        RECT 79.980 42.915 80.150 43.085 ;
        RECT 80.340 42.915 80.510 43.085 ;
        RECT 80.700 42.915 80.870 43.085 ;
        RECT 81.060 42.915 81.230 43.085 ;
        RECT 81.420 42.915 81.590 43.085 ;
        RECT 81.780 42.915 81.950 43.085 ;
        RECT 82.140 42.915 82.310 43.085 ;
        RECT 82.500 42.915 82.670 43.085 ;
        RECT 82.860 42.915 83.030 43.085 ;
        RECT 83.220 42.915 83.390 43.085 ;
        RECT 83.580 42.915 83.750 43.085 ;
        RECT 83.940 42.915 84.110 43.085 ;
        RECT 84.300 42.915 84.470 43.085 ;
        RECT 84.660 42.915 84.830 43.085 ;
        RECT 85.020 42.915 85.190 43.085 ;
        RECT 85.380 42.915 85.550 43.085 ;
        RECT 85.740 42.915 85.910 43.085 ;
        RECT 86.100 42.915 86.270 43.085 ;
        RECT 86.460 42.915 86.630 43.085 ;
        RECT 86.820 42.915 86.990 43.085 ;
        RECT 87.180 42.915 87.350 43.085 ;
        RECT 87.540 42.915 87.710 43.085 ;
        RECT 87.900 42.915 88.070 43.085 ;
        RECT 88.260 42.915 88.430 43.085 ;
        RECT 88.620 42.915 88.790 43.085 ;
        RECT 88.980 42.915 89.150 43.085 ;
        RECT 89.340 42.915 89.510 43.085 ;
        RECT 94.140 45.275 94.310 45.445 ;
        RECT 94.140 44.915 94.310 45.085 ;
        RECT 94.140 44.555 94.310 44.725 ;
        RECT 94.810 45.070 94.980 45.240 ;
        RECT 94.810 44.710 94.980 44.880 ;
        RECT 97.090 45.070 97.260 45.240 ;
        RECT 97.090 44.710 97.260 44.880 ;
        RECT 99.370 45.070 99.540 45.240 ;
        RECT 99.370 44.710 99.540 44.880 ;
        RECT 101.650 45.070 101.820 45.240 ;
        RECT 101.650 44.710 101.820 44.880 ;
        RECT 103.930 45.070 104.100 45.240 ;
        RECT 103.930 44.710 104.100 44.880 ;
        RECT 106.210 45.070 106.380 45.240 ;
        RECT 106.210 44.710 106.380 44.880 ;
        RECT 108.490 45.070 108.660 45.240 ;
        RECT 108.490 44.710 108.660 44.880 ;
        RECT 110.770 45.070 110.940 45.240 ;
        RECT 110.770 44.710 110.940 44.880 ;
        RECT 113.050 45.070 113.220 45.240 ;
        RECT 113.050 44.710 113.220 44.880 ;
        RECT 115.330 45.070 115.500 45.240 ;
        RECT 115.330 44.710 115.500 44.880 ;
        RECT 117.610 45.070 117.780 45.240 ;
        RECT 117.610 44.710 117.780 44.880 ;
        RECT 118.280 45.275 118.450 45.445 ;
        RECT 118.280 44.915 118.450 45.085 ;
        RECT 118.280 44.555 118.450 44.725 ;
        RECT 94.140 44.195 94.310 44.365 ;
        RECT 94.140 43.835 94.310 44.005 ;
        RECT 95.230 44.055 95.400 44.225 ;
        RECT 95.590 44.055 95.760 44.225 ;
        RECT 95.950 44.055 96.120 44.225 ;
        RECT 96.310 44.055 96.480 44.225 ;
        RECT 96.670 44.055 96.840 44.225 ;
        RECT 97.510 44.055 97.680 44.225 ;
        RECT 97.870 44.055 98.040 44.225 ;
        RECT 98.230 44.055 98.400 44.225 ;
        RECT 98.590 44.055 98.760 44.225 ;
        RECT 98.950 44.055 99.120 44.225 ;
        RECT 99.790 44.055 99.960 44.225 ;
        RECT 100.150 44.055 100.320 44.225 ;
        RECT 100.510 44.055 100.680 44.225 ;
        RECT 100.870 44.055 101.040 44.225 ;
        RECT 101.230 44.055 101.400 44.225 ;
        RECT 102.070 44.055 102.240 44.225 ;
        RECT 102.430 44.055 102.600 44.225 ;
        RECT 102.790 44.055 102.960 44.225 ;
        RECT 103.150 44.055 103.320 44.225 ;
        RECT 103.510 44.055 103.680 44.225 ;
        RECT 104.350 44.055 104.520 44.225 ;
        RECT 104.710 44.055 104.880 44.225 ;
        RECT 105.070 44.055 105.240 44.225 ;
        RECT 105.430 44.055 105.600 44.225 ;
        RECT 105.790 44.055 105.960 44.225 ;
        RECT 106.630 44.055 106.800 44.225 ;
        RECT 106.990 44.055 107.160 44.225 ;
        RECT 107.350 44.055 107.520 44.225 ;
        RECT 107.710 44.055 107.880 44.225 ;
        RECT 108.070 44.055 108.240 44.225 ;
        RECT 108.910 44.055 109.080 44.225 ;
        RECT 109.270 44.055 109.440 44.225 ;
        RECT 109.630 44.055 109.800 44.225 ;
        RECT 109.990 44.055 110.160 44.225 ;
        RECT 110.350 44.055 110.520 44.225 ;
        RECT 111.190 44.055 111.360 44.225 ;
        RECT 111.550 44.055 111.720 44.225 ;
        RECT 111.910 44.055 112.080 44.225 ;
        RECT 112.270 44.055 112.440 44.225 ;
        RECT 112.630 44.055 112.800 44.225 ;
        RECT 113.470 44.055 113.640 44.225 ;
        RECT 113.830 44.055 114.000 44.225 ;
        RECT 114.190 44.055 114.360 44.225 ;
        RECT 114.550 44.055 114.720 44.225 ;
        RECT 114.910 44.055 115.080 44.225 ;
        RECT 115.750 44.055 115.920 44.225 ;
        RECT 116.110 44.055 116.280 44.225 ;
        RECT 116.470 44.055 116.640 44.225 ;
        RECT 116.830 44.055 117.000 44.225 ;
        RECT 117.190 44.055 117.360 44.225 ;
        RECT 118.280 44.195 118.450 44.365 ;
        RECT 94.140 43.475 94.310 43.645 ;
        RECT 94.140 43.115 94.310 43.285 ;
        RECT 118.280 43.835 118.450 44.005 ;
        RECT 118.280 43.475 118.450 43.645 ;
        RECT 118.280 43.115 118.450 43.285 ;
        RECT 124.810 45.920 124.980 46.090 ;
        RECT 125.170 45.920 125.340 46.090 ;
        RECT 125.530 45.920 125.700 46.090 ;
        RECT 125.890 45.920 126.060 46.090 ;
        RECT 126.250 45.920 126.420 46.090 ;
        RECT 126.610 45.920 126.780 46.090 ;
        RECT 126.970 45.920 127.140 46.090 ;
        RECT 127.330 45.920 127.500 46.090 ;
        RECT 127.690 45.920 127.860 46.090 ;
        RECT 128.050 45.920 128.220 46.090 ;
        RECT 128.410 45.920 128.580 46.090 ;
        RECT 128.770 45.920 128.940 46.090 ;
        RECT 124.460 45.620 124.630 45.790 ;
        RECT 129.240 45.620 129.410 45.790 ;
        RECT 124.460 45.260 124.630 45.430 ;
        RECT 124.460 44.900 124.630 45.070 ;
        RECT 124.460 44.540 124.630 44.710 ;
        RECT 124.460 44.180 124.630 44.350 ;
        RECT 124.460 43.820 124.630 43.990 ;
        RECT 124.460 43.460 124.630 43.630 ;
        RECT 125.130 45.095 125.300 45.265 ;
        RECT 125.130 44.735 125.300 44.905 ;
        RECT 125.130 44.375 125.300 44.545 ;
        RECT 125.130 44.015 125.300 44.185 ;
        RECT 125.130 43.655 125.300 43.825 ;
        RECT 125.560 45.095 125.730 45.265 ;
        RECT 125.560 44.735 125.730 44.905 ;
        RECT 125.560 44.375 125.730 44.545 ;
        RECT 125.560 44.015 125.730 44.185 ;
        RECT 125.560 43.655 125.730 43.825 ;
        RECT 125.990 45.095 126.160 45.265 ;
        RECT 125.990 44.735 126.160 44.905 ;
        RECT 125.990 44.375 126.160 44.545 ;
        RECT 125.990 44.015 126.160 44.185 ;
        RECT 125.990 43.655 126.160 43.825 ;
        RECT 126.420 45.095 126.590 45.265 ;
        RECT 126.420 44.735 126.590 44.905 ;
        RECT 126.420 44.375 126.590 44.545 ;
        RECT 126.420 44.015 126.590 44.185 ;
        RECT 126.420 43.655 126.590 43.825 ;
        RECT 126.850 45.095 127.020 45.265 ;
        RECT 126.850 44.735 127.020 44.905 ;
        RECT 126.850 44.375 127.020 44.545 ;
        RECT 126.850 44.015 127.020 44.185 ;
        RECT 126.850 43.655 127.020 43.825 ;
        RECT 127.280 45.095 127.450 45.265 ;
        RECT 127.280 44.735 127.450 44.905 ;
        RECT 127.280 44.375 127.450 44.545 ;
        RECT 127.280 44.015 127.450 44.185 ;
        RECT 127.280 43.655 127.450 43.825 ;
        RECT 127.710 45.095 127.880 45.265 ;
        RECT 127.710 44.735 127.880 44.905 ;
        RECT 127.710 44.375 127.880 44.545 ;
        RECT 127.710 44.015 127.880 44.185 ;
        RECT 127.710 43.655 127.880 43.825 ;
        RECT 128.140 45.095 128.310 45.265 ;
        RECT 128.140 44.735 128.310 44.905 ;
        RECT 128.140 44.375 128.310 44.545 ;
        RECT 128.140 44.015 128.310 44.185 ;
        RECT 128.140 43.655 128.310 43.825 ;
        RECT 128.570 45.095 128.740 45.265 ;
        RECT 128.570 44.735 128.740 44.905 ;
        RECT 128.570 44.375 128.740 44.545 ;
        RECT 128.570 44.015 128.740 44.185 ;
        RECT 128.570 43.655 128.740 43.825 ;
        RECT 129.240 45.260 129.410 45.430 ;
        RECT 129.240 44.900 129.410 45.070 ;
        RECT 129.240 44.540 129.410 44.710 ;
        RECT 129.240 44.180 129.410 44.350 ;
        RECT 129.240 43.820 129.410 43.990 ;
        RECT 129.240 43.460 129.410 43.630 ;
        RECT 124.460 43.100 124.630 43.270 ;
        RECT 125.380 43.040 125.550 43.210 ;
        RECT 125.740 43.040 125.910 43.210 ;
        RECT 126.240 43.040 126.410 43.210 ;
        RECT 126.600 43.040 126.770 43.210 ;
        RECT 127.100 43.040 127.270 43.210 ;
        RECT 127.460 43.040 127.630 43.210 ;
        RECT 127.960 43.040 128.130 43.210 ;
        RECT 128.320 43.040 128.490 43.210 ;
        RECT 129.240 43.100 129.410 43.270 ;
        RECT 135.470 45.920 135.640 46.090 ;
        RECT 135.830 45.920 136.000 46.090 ;
        RECT 136.190 45.920 136.360 46.090 ;
        RECT 136.550 45.920 136.720 46.090 ;
        RECT 136.910 45.920 137.080 46.090 ;
        RECT 137.270 45.920 137.440 46.090 ;
        RECT 137.630 45.920 137.800 46.090 ;
        RECT 137.990 45.920 138.160 46.090 ;
        RECT 138.350 45.920 138.520 46.090 ;
        RECT 138.710 45.920 138.880 46.090 ;
        RECT 139.070 45.920 139.240 46.090 ;
        RECT 139.430 45.920 139.600 46.090 ;
        RECT 139.790 45.920 139.960 46.090 ;
        RECT 140.150 45.920 140.320 46.090 ;
        RECT 140.510 45.920 140.680 46.090 ;
        RECT 140.870 45.920 141.040 46.090 ;
        RECT 141.230 45.920 141.400 46.090 ;
        RECT 141.590 45.920 141.760 46.090 ;
        RECT 141.950 45.920 142.120 46.090 ;
        RECT 142.310 45.920 142.480 46.090 ;
        RECT 142.670 45.920 142.840 46.090 ;
        RECT 143.030 45.920 143.200 46.090 ;
        RECT 143.390 45.920 143.560 46.090 ;
        RECT 143.750 45.920 143.920 46.090 ;
        RECT 135.120 45.620 135.290 45.790 ;
        RECT 144.200 45.620 144.370 45.790 ;
        RECT 135.120 45.260 135.290 45.430 ;
        RECT 135.120 44.900 135.290 45.070 ;
        RECT 135.120 44.540 135.290 44.710 ;
        RECT 135.120 44.180 135.290 44.350 ;
        RECT 135.120 43.820 135.290 43.990 ;
        RECT 135.120 43.460 135.290 43.630 ;
        RECT 135.790 45.095 135.960 45.265 ;
        RECT 135.790 44.735 135.960 44.905 ;
        RECT 135.790 44.375 135.960 44.545 ;
        RECT 135.790 44.015 135.960 44.185 ;
        RECT 135.790 43.655 135.960 43.825 ;
        RECT 136.220 45.095 136.390 45.265 ;
        RECT 136.220 44.735 136.390 44.905 ;
        RECT 136.220 44.375 136.390 44.545 ;
        RECT 136.220 44.015 136.390 44.185 ;
        RECT 136.220 43.655 136.390 43.825 ;
        RECT 136.650 45.095 136.820 45.265 ;
        RECT 136.650 44.735 136.820 44.905 ;
        RECT 136.650 44.375 136.820 44.545 ;
        RECT 136.650 44.015 136.820 44.185 ;
        RECT 136.650 43.655 136.820 43.825 ;
        RECT 137.080 45.095 137.250 45.265 ;
        RECT 137.080 44.735 137.250 44.905 ;
        RECT 137.080 44.375 137.250 44.545 ;
        RECT 137.080 44.015 137.250 44.185 ;
        RECT 137.080 43.655 137.250 43.825 ;
        RECT 137.510 45.095 137.680 45.265 ;
        RECT 137.510 44.735 137.680 44.905 ;
        RECT 137.510 44.375 137.680 44.545 ;
        RECT 137.510 44.015 137.680 44.185 ;
        RECT 137.510 43.655 137.680 43.825 ;
        RECT 137.940 45.095 138.110 45.265 ;
        RECT 137.940 44.735 138.110 44.905 ;
        RECT 137.940 44.375 138.110 44.545 ;
        RECT 137.940 44.015 138.110 44.185 ;
        RECT 137.940 43.655 138.110 43.825 ;
        RECT 138.370 45.095 138.540 45.265 ;
        RECT 138.370 44.735 138.540 44.905 ;
        RECT 138.370 44.375 138.540 44.545 ;
        RECT 138.370 44.015 138.540 44.185 ;
        RECT 138.370 43.655 138.540 43.825 ;
        RECT 138.800 45.095 138.970 45.265 ;
        RECT 138.800 44.735 138.970 44.905 ;
        RECT 138.800 44.375 138.970 44.545 ;
        RECT 138.800 44.015 138.970 44.185 ;
        RECT 138.800 43.655 138.970 43.825 ;
        RECT 139.230 45.095 139.400 45.265 ;
        RECT 139.230 44.735 139.400 44.905 ;
        RECT 139.230 44.375 139.400 44.545 ;
        RECT 139.230 44.015 139.400 44.185 ;
        RECT 139.230 43.655 139.400 43.825 ;
        RECT 139.660 45.095 139.830 45.265 ;
        RECT 139.660 44.735 139.830 44.905 ;
        RECT 139.660 44.375 139.830 44.545 ;
        RECT 139.660 44.015 139.830 44.185 ;
        RECT 139.660 43.655 139.830 43.825 ;
        RECT 140.090 45.095 140.260 45.265 ;
        RECT 140.090 44.735 140.260 44.905 ;
        RECT 140.090 44.375 140.260 44.545 ;
        RECT 140.090 44.015 140.260 44.185 ;
        RECT 140.090 43.655 140.260 43.825 ;
        RECT 140.520 45.095 140.690 45.265 ;
        RECT 140.520 44.735 140.690 44.905 ;
        RECT 140.520 44.375 140.690 44.545 ;
        RECT 140.520 44.015 140.690 44.185 ;
        RECT 140.520 43.655 140.690 43.825 ;
        RECT 140.950 45.095 141.120 45.265 ;
        RECT 140.950 44.735 141.120 44.905 ;
        RECT 140.950 44.375 141.120 44.545 ;
        RECT 140.950 44.015 141.120 44.185 ;
        RECT 140.950 43.655 141.120 43.825 ;
        RECT 141.380 45.095 141.550 45.265 ;
        RECT 141.380 44.735 141.550 44.905 ;
        RECT 141.380 44.375 141.550 44.545 ;
        RECT 141.380 44.015 141.550 44.185 ;
        RECT 141.380 43.655 141.550 43.825 ;
        RECT 141.810 45.095 141.980 45.265 ;
        RECT 141.810 44.735 141.980 44.905 ;
        RECT 141.810 44.375 141.980 44.545 ;
        RECT 141.810 44.015 141.980 44.185 ;
        RECT 141.810 43.655 141.980 43.825 ;
        RECT 142.240 45.095 142.410 45.265 ;
        RECT 142.240 44.735 142.410 44.905 ;
        RECT 142.240 44.375 142.410 44.545 ;
        RECT 142.240 44.015 142.410 44.185 ;
        RECT 142.240 43.655 142.410 43.825 ;
        RECT 142.670 45.095 142.840 45.265 ;
        RECT 142.670 44.735 142.840 44.905 ;
        RECT 142.670 44.375 142.840 44.545 ;
        RECT 142.670 44.015 142.840 44.185 ;
        RECT 142.670 43.655 142.840 43.825 ;
        RECT 143.100 45.095 143.270 45.265 ;
        RECT 143.100 44.735 143.270 44.905 ;
        RECT 143.100 44.375 143.270 44.545 ;
        RECT 143.100 44.015 143.270 44.185 ;
        RECT 143.100 43.655 143.270 43.825 ;
        RECT 143.530 45.095 143.700 45.265 ;
        RECT 143.530 44.735 143.700 44.905 ;
        RECT 143.530 44.375 143.700 44.545 ;
        RECT 143.530 44.015 143.700 44.185 ;
        RECT 143.530 43.655 143.700 43.825 ;
        RECT 144.200 45.260 144.370 45.430 ;
        RECT 144.200 44.900 144.370 45.070 ;
        RECT 144.200 44.540 144.370 44.710 ;
        RECT 144.200 44.180 144.370 44.350 ;
        RECT 144.200 43.820 144.370 43.990 ;
        RECT 144.200 43.460 144.370 43.630 ;
        RECT 135.120 43.100 135.290 43.270 ;
        RECT 136.040 43.040 136.210 43.210 ;
        RECT 136.400 43.040 136.570 43.210 ;
        RECT 136.900 43.040 137.070 43.210 ;
        RECT 137.260 43.040 137.430 43.210 ;
        RECT 137.760 43.040 137.930 43.210 ;
        RECT 138.120 43.040 138.290 43.210 ;
        RECT 138.620 43.040 138.790 43.210 ;
        RECT 138.980 43.040 139.150 43.210 ;
        RECT 139.480 43.040 139.650 43.210 ;
        RECT 139.840 43.040 140.010 43.210 ;
        RECT 140.340 43.040 140.510 43.210 ;
        RECT 140.700 43.040 140.870 43.210 ;
        RECT 141.200 43.040 141.370 43.210 ;
        RECT 141.560 43.040 141.730 43.210 ;
        RECT 142.060 43.040 142.230 43.210 ;
        RECT 142.420 43.040 142.590 43.210 ;
        RECT 142.920 43.040 143.090 43.210 ;
        RECT 143.280 43.040 143.450 43.210 ;
        RECT 144.200 43.100 144.370 43.270 ;
        RECT 94.140 41.645 94.310 41.815 ;
        RECT 69.540 41.430 69.710 41.600 ;
        RECT 69.900 41.430 70.070 41.600 ;
        RECT 70.260 41.430 70.430 41.600 ;
        RECT 70.620 41.430 70.790 41.600 ;
        RECT 70.980 41.430 71.150 41.600 ;
        RECT 71.340 41.430 71.510 41.600 ;
        RECT 71.700 41.430 71.870 41.600 ;
        RECT 72.060 41.430 72.230 41.600 ;
        RECT 72.420 41.430 72.590 41.600 ;
        RECT 72.780 41.430 72.950 41.600 ;
        RECT 73.140 41.430 73.310 41.600 ;
        RECT 73.500 41.430 73.670 41.600 ;
        RECT 73.860 41.430 74.030 41.600 ;
        RECT 74.220 41.430 74.390 41.600 ;
        RECT 74.580 41.430 74.750 41.600 ;
        RECT 74.940 41.430 75.110 41.600 ;
        RECT 75.300 41.430 75.470 41.600 ;
        RECT 75.660 41.430 75.830 41.600 ;
        RECT 76.020 41.430 76.190 41.600 ;
        RECT 76.380 41.430 76.550 41.600 ;
        RECT 76.740 41.430 76.910 41.600 ;
        RECT 77.100 41.430 77.270 41.600 ;
        RECT 77.460 41.430 77.630 41.600 ;
        RECT 77.820 41.430 77.990 41.600 ;
        RECT 78.180 41.430 78.350 41.600 ;
        RECT 78.540 41.430 78.710 41.600 ;
        RECT 78.900 41.430 79.070 41.600 ;
        RECT 79.260 41.430 79.430 41.600 ;
        RECT 79.620 41.430 79.790 41.600 ;
        RECT 79.980 41.430 80.150 41.600 ;
        RECT 80.340 41.430 80.510 41.600 ;
        RECT 80.700 41.430 80.870 41.600 ;
        RECT 81.060 41.430 81.230 41.600 ;
        RECT 81.420 41.430 81.590 41.600 ;
        RECT 81.780 41.430 81.950 41.600 ;
        RECT 82.140 41.430 82.310 41.600 ;
        RECT 82.500 41.430 82.670 41.600 ;
        RECT 82.860 41.430 83.030 41.600 ;
        RECT 83.220 41.430 83.390 41.600 ;
        RECT 83.580 41.430 83.750 41.600 ;
        RECT 83.940 41.430 84.110 41.600 ;
        RECT 84.300 41.430 84.470 41.600 ;
        RECT 84.660 41.430 84.830 41.600 ;
        RECT 85.020 41.430 85.190 41.600 ;
        RECT 85.380 41.430 85.550 41.600 ;
        RECT 85.740 41.430 85.910 41.600 ;
        RECT 86.100 41.430 86.270 41.600 ;
        RECT 86.460 41.430 86.630 41.600 ;
        RECT 86.820 41.430 86.990 41.600 ;
        RECT 87.180 41.430 87.350 41.600 ;
        RECT 87.540 41.430 87.710 41.600 ;
        RECT 87.900 41.430 88.070 41.600 ;
        RECT 88.260 41.430 88.430 41.600 ;
        RECT 88.620 41.430 88.790 41.600 ;
        RECT 88.980 41.430 89.150 41.600 ;
        RECT 89.340 41.430 89.510 41.600 ;
        RECT 69.190 41.120 69.360 41.290 ;
        RECT 69.190 40.760 69.360 40.930 ;
        RECT 70.245 40.880 70.415 41.050 ;
        RECT 70.605 40.880 70.775 41.050 ;
        RECT 70.965 40.880 71.135 41.050 ;
        RECT 71.325 40.880 71.495 41.050 ;
        RECT 71.685 40.880 71.855 41.050 ;
        RECT 72.045 40.880 72.215 41.050 ;
        RECT 72.840 40.880 73.010 41.050 ;
        RECT 73.200 40.880 73.370 41.050 ;
        RECT 73.560 40.880 73.730 41.050 ;
        RECT 73.920 40.880 74.090 41.050 ;
        RECT 74.280 40.880 74.450 41.050 ;
        RECT 75.120 40.880 75.290 41.050 ;
        RECT 75.480 40.880 75.650 41.050 ;
        RECT 75.840 40.880 76.010 41.050 ;
        RECT 76.200 40.880 76.370 41.050 ;
        RECT 76.560 40.880 76.730 41.050 ;
        RECT 77.365 40.880 77.535 41.050 ;
        RECT 77.725 40.880 77.895 41.050 ;
        RECT 78.085 40.880 78.255 41.050 ;
        RECT 78.445 40.880 78.615 41.050 ;
        RECT 78.805 40.880 78.975 41.050 ;
        RECT 79.165 40.880 79.335 41.050 ;
        RECT 79.925 40.880 80.095 41.050 ;
        RECT 80.285 40.880 80.455 41.050 ;
        RECT 80.645 40.880 80.815 41.050 ;
        RECT 81.005 40.880 81.175 41.050 ;
        RECT 81.365 40.880 81.535 41.050 ;
        RECT 81.725 40.880 81.895 41.050 ;
        RECT 87.045 40.880 87.215 41.050 ;
        RECT 87.405 40.880 87.575 41.050 ;
        RECT 87.765 40.880 87.935 41.050 ;
        RECT 88.125 40.880 88.295 41.050 ;
        RECT 88.485 40.880 88.655 41.050 ;
        RECT 88.845 40.880 89.015 41.050 ;
        RECT 89.890 41.120 90.060 41.290 ;
        RECT 89.890 40.760 90.060 40.930 ;
        RECT 69.190 40.400 69.360 40.570 ;
        RECT 69.190 40.040 69.360 40.210 ;
        RECT 69.190 39.680 69.360 39.850 ;
        RECT 69.860 40.225 70.030 40.395 ;
        RECT 69.860 39.865 70.030 40.035 ;
        RECT 71.140 40.225 71.310 40.395 ;
        RECT 71.140 39.865 71.310 40.035 ;
        RECT 72.420 40.225 72.590 40.395 ;
        RECT 72.420 39.865 72.590 40.035 ;
        RECT 74.700 40.225 74.870 40.395 ;
        RECT 74.700 39.865 74.870 40.035 ;
        RECT 76.980 40.225 77.150 40.395 ;
        RECT 76.980 39.865 77.150 40.035 ;
        RECT 78.260 40.225 78.430 40.395 ;
        RECT 78.260 39.865 78.430 40.035 ;
        RECT 79.540 40.225 79.710 40.395 ;
        RECT 79.540 39.865 79.710 40.035 ;
        RECT 80.820 40.225 80.990 40.395 ;
        RECT 80.820 39.865 80.990 40.035 ;
        RECT 82.100 40.225 82.270 40.395 ;
        RECT 82.100 39.865 82.270 40.035 ;
        RECT 84.380 40.225 84.550 40.395 ;
        RECT 84.380 39.865 84.550 40.035 ;
        RECT 86.660 40.225 86.830 40.395 ;
        RECT 86.660 39.865 86.830 40.035 ;
        RECT 87.940 40.225 88.110 40.395 ;
        RECT 87.940 39.865 88.110 40.035 ;
        RECT 89.220 40.225 89.390 40.395 ;
        RECT 89.220 39.865 89.390 40.035 ;
        RECT 89.890 40.400 90.060 40.570 ;
        RECT 89.890 40.040 90.060 40.210 ;
        RECT 89.890 39.680 90.060 39.850 ;
        RECT 69.190 39.320 69.360 39.490 ;
        RECT 94.140 41.285 94.310 41.455 ;
        RECT 118.280 41.645 118.450 41.815 ;
        RECT 118.280 41.285 118.450 41.455 ;
        RECT 94.140 40.925 94.310 41.095 ;
        RECT 95.230 40.925 95.400 41.095 ;
        RECT 95.590 40.925 95.760 41.095 ;
        RECT 95.950 40.925 96.120 41.095 ;
        RECT 96.310 40.925 96.480 41.095 ;
        RECT 96.670 40.925 96.840 41.095 ;
        RECT 97.510 40.925 97.680 41.095 ;
        RECT 97.870 40.925 98.040 41.095 ;
        RECT 98.230 40.925 98.400 41.095 ;
        RECT 98.590 40.925 98.760 41.095 ;
        RECT 98.950 40.925 99.120 41.095 ;
        RECT 99.790 40.925 99.960 41.095 ;
        RECT 100.150 40.925 100.320 41.095 ;
        RECT 100.510 40.925 100.680 41.095 ;
        RECT 100.870 40.925 101.040 41.095 ;
        RECT 101.230 40.925 101.400 41.095 ;
        RECT 102.070 40.925 102.240 41.095 ;
        RECT 102.430 40.925 102.600 41.095 ;
        RECT 102.790 40.925 102.960 41.095 ;
        RECT 103.150 40.925 103.320 41.095 ;
        RECT 103.510 40.925 103.680 41.095 ;
        RECT 104.350 40.925 104.520 41.095 ;
        RECT 104.710 40.925 104.880 41.095 ;
        RECT 105.070 40.925 105.240 41.095 ;
        RECT 105.430 40.925 105.600 41.095 ;
        RECT 105.790 40.925 105.960 41.095 ;
        RECT 106.630 40.925 106.800 41.095 ;
        RECT 106.990 40.925 107.160 41.095 ;
        RECT 107.350 40.925 107.520 41.095 ;
        RECT 107.710 40.925 107.880 41.095 ;
        RECT 108.070 40.925 108.240 41.095 ;
        RECT 108.910 40.925 109.080 41.095 ;
        RECT 109.270 40.925 109.440 41.095 ;
        RECT 109.630 40.925 109.800 41.095 ;
        RECT 109.990 40.925 110.160 41.095 ;
        RECT 110.350 40.925 110.520 41.095 ;
        RECT 111.190 40.925 111.360 41.095 ;
        RECT 111.550 40.925 111.720 41.095 ;
        RECT 111.910 40.925 112.080 41.095 ;
        RECT 112.270 40.925 112.440 41.095 ;
        RECT 112.630 40.925 112.800 41.095 ;
        RECT 113.470 40.925 113.640 41.095 ;
        RECT 113.830 40.925 114.000 41.095 ;
        RECT 114.190 40.925 114.360 41.095 ;
        RECT 114.550 40.925 114.720 41.095 ;
        RECT 114.910 40.925 115.080 41.095 ;
        RECT 115.750 40.925 115.920 41.095 ;
        RECT 116.110 40.925 116.280 41.095 ;
        RECT 116.470 40.925 116.640 41.095 ;
        RECT 116.830 40.925 117.000 41.095 ;
        RECT 117.190 40.925 117.360 41.095 ;
        RECT 118.280 40.925 118.450 41.095 ;
        RECT 94.140 40.565 94.310 40.735 ;
        RECT 94.140 40.205 94.310 40.375 ;
        RECT 94.810 40.340 94.980 40.510 ;
        RECT 97.090 40.340 97.260 40.510 ;
        RECT 99.370 40.340 99.540 40.510 ;
        RECT 101.650 40.340 101.820 40.510 ;
        RECT 103.930 40.340 104.100 40.510 ;
        RECT 106.210 40.340 106.380 40.510 ;
        RECT 108.490 40.340 108.660 40.510 ;
        RECT 110.770 40.340 110.940 40.510 ;
        RECT 113.050 40.340 113.220 40.510 ;
        RECT 115.330 40.340 115.500 40.510 ;
        RECT 117.610 40.340 117.780 40.510 ;
        RECT 118.280 40.565 118.450 40.735 ;
        RECT 118.280 40.205 118.450 40.375 ;
        RECT 94.140 39.845 94.310 40.015 ;
        RECT 118.280 39.845 118.450 40.015 ;
        RECT 94.490 39.545 94.660 39.715 ;
        RECT 94.850 39.545 95.020 39.715 ;
        RECT 95.210 39.545 95.380 39.715 ;
        RECT 95.570 39.545 95.740 39.715 ;
        RECT 95.930 39.545 96.100 39.715 ;
        RECT 96.290 39.545 96.460 39.715 ;
        RECT 96.650 39.545 96.820 39.715 ;
        RECT 97.010 39.545 97.180 39.715 ;
        RECT 97.370 39.545 97.540 39.715 ;
        RECT 97.730 39.545 97.900 39.715 ;
        RECT 98.090 39.545 98.260 39.715 ;
        RECT 98.450 39.545 98.620 39.715 ;
        RECT 98.810 39.545 98.980 39.715 ;
        RECT 99.170 39.545 99.340 39.715 ;
        RECT 99.530 39.545 99.700 39.715 ;
        RECT 99.890 39.545 100.060 39.715 ;
        RECT 100.250 39.545 100.420 39.715 ;
        RECT 100.610 39.545 100.780 39.715 ;
        RECT 100.970 39.545 101.140 39.715 ;
        RECT 101.330 39.545 101.500 39.715 ;
        RECT 101.690 39.545 101.860 39.715 ;
        RECT 102.050 39.545 102.220 39.715 ;
        RECT 102.410 39.545 102.580 39.715 ;
        RECT 102.770 39.545 102.940 39.715 ;
        RECT 103.130 39.545 103.300 39.715 ;
        RECT 103.490 39.545 103.660 39.715 ;
        RECT 103.850 39.545 104.020 39.715 ;
        RECT 104.210 39.545 104.380 39.715 ;
        RECT 104.570 39.545 104.740 39.715 ;
        RECT 104.930 39.545 105.100 39.715 ;
        RECT 105.290 39.545 105.460 39.715 ;
        RECT 105.650 39.545 105.820 39.715 ;
        RECT 106.010 39.545 106.180 39.715 ;
        RECT 106.370 39.545 106.540 39.715 ;
        RECT 106.730 39.545 106.900 39.715 ;
        RECT 107.090 39.545 107.260 39.715 ;
        RECT 107.450 39.545 107.620 39.715 ;
        RECT 107.810 39.545 107.980 39.715 ;
        RECT 108.170 39.545 108.340 39.715 ;
        RECT 108.530 39.545 108.700 39.715 ;
        RECT 108.890 39.545 109.060 39.715 ;
        RECT 109.250 39.545 109.420 39.715 ;
        RECT 109.610 39.545 109.780 39.715 ;
        RECT 109.970 39.545 110.140 39.715 ;
        RECT 110.330 39.545 110.500 39.715 ;
        RECT 110.690 39.545 110.860 39.715 ;
        RECT 111.050 39.545 111.220 39.715 ;
        RECT 111.410 39.545 111.580 39.715 ;
        RECT 111.770 39.545 111.940 39.715 ;
        RECT 112.130 39.545 112.300 39.715 ;
        RECT 112.490 39.545 112.660 39.715 ;
        RECT 112.850 39.545 113.020 39.715 ;
        RECT 113.210 39.545 113.380 39.715 ;
        RECT 113.570 39.545 113.740 39.715 ;
        RECT 113.930 39.545 114.100 39.715 ;
        RECT 114.290 39.545 114.460 39.715 ;
        RECT 114.650 39.545 114.820 39.715 ;
        RECT 115.010 39.545 115.180 39.715 ;
        RECT 115.370 39.545 115.540 39.715 ;
        RECT 115.730 39.545 115.900 39.715 ;
        RECT 116.090 39.545 116.260 39.715 ;
        RECT 116.450 39.545 116.620 39.715 ;
        RECT 116.810 39.545 116.980 39.715 ;
        RECT 117.170 39.545 117.340 39.715 ;
        RECT 117.530 39.545 117.700 39.715 ;
        RECT 117.890 39.545 118.060 39.715 ;
        RECT 124.460 41.605 124.630 41.775 ;
        RECT 124.460 41.245 124.630 41.415 ;
        RECT 125.380 41.360 125.550 41.530 ;
        RECT 125.740 41.360 125.910 41.530 ;
        RECT 126.240 41.360 126.410 41.530 ;
        RECT 126.600 41.360 126.770 41.530 ;
        RECT 127.100 41.360 127.270 41.530 ;
        RECT 127.460 41.360 127.630 41.530 ;
        RECT 127.960 41.360 128.130 41.530 ;
        RECT 128.320 41.360 128.490 41.530 ;
        RECT 129.240 41.605 129.410 41.775 ;
        RECT 129.240 41.245 129.410 41.415 ;
        RECT 124.460 40.885 124.630 41.055 ;
        RECT 124.460 40.525 124.630 40.695 ;
        RECT 124.460 40.165 124.630 40.335 ;
        RECT 125.130 40.705 125.300 40.875 ;
        RECT 125.130 40.345 125.300 40.515 ;
        RECT 125.560 40.705 125.730 40.875 ;
        RECT 125.560 40.345 125.730 40.515 ;
        RECT 125.990 40.705 126.160 40.875 ;
        RECT 125.990 40.345 126.160 40.515 ;
        RECT 126.420 40.705 126.590 40.875 ;
        RECT 126.420 40.345 126.590 40.515 ;
        RECT 126.850 40.705 127.020 40.875 ;
        RECT 126.850 40.345 127.020 40.515 ;
        RECT 127.280 40.705 127.450 40.875 ;
        RECT 127.280 40.345 127.450 40.515 ;
        RECT 127.710 40.705 127.880 40.875 ;
        RECT 127.710 40.345 127.880 40.515 ;
        RECT 128.140 40.705 128.310 40.875 ;
        RECT 128.140 40.345 128.310 40.515 ;
        RECT 128.570 40.705 128.740 40.875 ;
        RECT 128.570 40.345 128.740 40.515 ;
        RECT 129.240 40.885 129.410 41.055 ;
        RECT 129.240 40.525 129.410 40.695 ;
        RECT 129.240 40.165 129.410 40.335 ;
        RECT 124.460 39.805 124.630 39.975 ;
        RECT 129.240 39.805 129.410 39.975 ;
        RECT 124.810 39.505 124.980 39.675 ;
        RECT 125.170 39.505 125.340 39.675 ;
        RECT 125.530 39.505 125.700 39.675 ;
        RECT 125.890 39.505 126.060 39.675 ;
        RECT 126.250 39.505 126.420 39.675 ;
        RECT 126.610 39.505 126.780 39.675 ;
        RECT 126.970 39.505 127.140 39.675 ;
        RECT 127.330 39.505 127.500 39.675 ;
        RECT 127.690 39.505 127.860 39.675 ;
        RECT 128.050 39.505 128.220 39.675 ;
        RECT 128.410 39.505 128.580 39.675 ;
        RECT 128.770 39.505 128.940 39.675 ;
        RECT 135.120 41.605 135.290 41.775 ;
        RECT 135.120 41.245 135.290 41.415 ;
        RECT 136.040 41.360 136.210 41.530 ;
        RECT 136.400 41.360 136.570 41.530 ;
        RECT 136.900 41.360 137.070 41.530 ;
        RECT 137.260 41.360 137.430 41.530 ;
        RECT 137.760 41.360 137.930 41.530 ;
        RECT 138.120 41.360 138.290 41.530 ;
        RECT 138.620 41.360 138.790 41.530 ;
        RECT 138.980 41.360 139.150 41.530 ;
        RECT 139.480 41.360 139.650 41.530 ;
        RECT 139.840 41.360 140.010 41.530 ;
        RECT 140.340 41.360 140.510 41.530 ;
        RECT 140.700 41.360 140.870 41.530 ;
        RECT 141.200 41.360 141.370 41.530 ;
        RECT 141.560 41.360 141.730 41.530 ;
        RECT 142.060 41.360 142.230 41.530 ;
        RECT 142.420 41.360 142.590 41.530 ;
        RECT 142.920 41.360 143.090 41.530 ;
        RECT 143.280 41.360 143.450 41.530 ;
        RECT 144.200 41.605 144.370 41.775 ;
        RECT 144.200 41.245 144.370 41.415 ;
        RECT 135.120 40.885 135.290 41.055 ;
        RECT 135.120 40.525 135.290 40.695 ;
        RECT 135.120 40.165 135.290 40.335 ;
        RECT 135.790 40.705 135.960 40.875 ;
        RECT 135.790 40.345 135.960 40.515 ;
        RECT 136.220 40.705 136.390 40.875 ;
        RECT 136.220 40.345 136.390 40.515 ;
        RECT 136.650 40.705 136.820 40.875 ;
        RECT 136.650 40.345 136.820 40.515 ;
        RECT 137.080 40.705 137.250 40.875 ;
        RECT 137.080 40.345 137.250 40.515 ;
        RECT 137.510 40.705 137.680 40.875 ;
        RECT 137.510 40.345 137.680 40.515 ;
        RECT 137.940 40.705 138.110 40.875 ;
        RECT 137.940 40.345 138.110 40.515 ;
        RECT 138.370 40.705 138.540 40.875 ;
        RECT 138.370 40.345 138.540 40.515 ;
        RECT 138.800 40.705 138.970 40.875 ;
        RECT 138.800 40.345 138.970 40.515 ;
        RECT 139.230 40.705 139.400 40.875 ;
        RECT 139.230 40.345 139.400 40.515 ;
        RECT 139.660 40.705 139.830 40.875 ;
        RECT 139.660 40.345 139.830 40.515 ;
        RECT 140.090 40.705 140.260 40.875 ;
        RECT 140.090 40.345 140.260 40.515 ;
        RECT 140.520 40.705 140.690 40.875 ;
        RECT 140.520 40.345 140.690 40.515 ;
        RECT 140.950 40.705 141.120 40.875 ;
        RECT 140.950 40.345 141.120 40.515 ;
        RECT 141.380 40.705 141.550 40.875 ;
        RECT 141.380 40.345 141.550 40.515 ;
        RECT 141.810 40.705 141.980 40.875 ;
        RECT 141.810 40.345 141.980 40.515 ;
        RECT 142.240 40.705 142.410 40.875 ;
        RECT 142.240 40.345 142.410 40.515 ;
        RECT 142.670 40.705 142.840 40.875 ;
        RECT 142.670 40.345 142.840 40.515 ;
        RECT 143.100 40.705 143.270 40.875 ;
        RECT 143.100 40.345 143.270 40.515 ;
        RECT 143.530 40.705 143.700 40.875 ;
        RECT 143.530 40.345 143.700 40.515 ;
        RECT 144.200 40.885 144.370 41.055 ;
        RECT 144.200 40.525 144.370 40.695 ;
        RECT 144.200 40.165 144.370 40.335 ;
        RECT 135.120 39.805 135.290 39.975 ;
        RECT 144.200 39.805 144.370 39.975 ;
        RECT 135.470 39.505 135.640 39.675 ;
        RECT 135.830 39.505 136.000 39.675 ;
        RECT 136.190 39.505 136.360 39.675 ;
        RECT 136.550 39.505 136.720 39.675 ;
        RECT 136.910 39.505 137.080 39.675 ;
        RECT 137.270 39.505 137.440 39.675 ;
        RECT 137.630 39.505 137.800 39.675 ;
        RECT 137.990 39.505 138.160 39.675 ;
        RECT 138.350 39.505 138.520 39.675 ;
        RECT 138.710 39.505 138.880 39.675 ;
        RECT 139.070 39.505 139.240 39.675 ;
        RECT 139.430 39.505 139.600 39.675 ;
        RECT 139.790 39.505 139.960 39.675 ;
        RECT 140.150 39.505 140.320 39.675 ;
        RECT 140.510 39.505 140.680 39.675 ;
        RECT 140.870 39.505 141.040 39.675 ;
        RECT 141.230 39.505 141.400 39.675 ;
        RECT 141.590 39.505 141.760 39.675 ;
        RECT 141.950 39.505 142.120 39.675 ;
        RECT 142.310 39.505 142.480 39.675 ;
        RECT 142.670 39.505 142.840 39.675 ;
        RECT 143.030 39.505 143.200 39.675 ;
        RECT 143.390 39.505 143.560 39.675 ;
        RECT 143.750 39.505 143.920 39.675 ;
        RECT 70.245 39.210 70.415 39.380 ;
        RECT 70.605 39.210 70.775 39.380 ;
        RECT 70.965 39.210 71.135 39.380 ;
        RECT 71.325 39.210 71.495 39.380 ;
        RECT 71.685 39.210 71.855 39.380 ;
        RECT 72.045 39.210 72.215 39.380 ;
        RECT 72.840 39.210 73.010 39.380 ;
        RECT 73.200 39.210 73.370 39.380 ;
        RECT 73.560 39.210 73.730 39.380 ;
        RECT 73.920 39.210 74.090 39.380 ;
        RECT 74.280 39.210 74.450 39.380 ;
        RECT 75.120 39.210 75.290 39.380 ;
        RECT 75.480 39.210 75.650 39.380 ;
        RECT 75.840 39.210 76.010 39.380 ;
        RECT 76.200 39.210 76.370 39.380 ;
        RECT 76.560 39.210 76.730 39.380 ;
        RECT 77.365 39.210 77.535 39.380 ;
        RECT 77.725 39.210 77.895 39.380 ;
        RECT 78.085 39.210 78.255 39.380 ;
        RECT 78.445 39.210 78.615 39.380 ;
        RECT 78.805 39.210 78.975 39.380 ;
        RECT 79.165 39.210 79.335 39.380 ;
        RECT 79.925 39.210 80.095 39.380 ;
        RECT 80.285 39.210 80.455 39.380 ;
        RECT 80.645 39.210 80.815 39.380 ;
        RECT 81.005 39.210 81.175 39.380 ;
        RECT 81.365 39.210 81.535 39.380 ;
        RECT 81.725 39.210 81.895 39.380 ;
        RECT 82.520 39.210 82.690 39.380 ;
        RECT 82.880 39.210 83.050 39.380 ;
        RECT 83.240 39.210 83.410 39.380 ;
        RECT 83.600 39.210 83.770 39.380 ;
        RECT 83.960 39.210 84.130 39.380 ;
        RECT 84.800 39.210 84.970 39.380 ;
        RECT 85.160 39.210 85.330 39.380 ;
        RECT 85.520 39.210 85.690 39.380 ;
        RECT 85.880 39.210 86.050 39.380 ;
        RECT 86.240 39.210 86.410 39.380 ;
        RECT 87.045 39.210 87.215 39.380 ;
        RECT 87.405 39.210 87.575 39.380 ;
        RECT 87.765 39.210 87.935 39.380 ;
        RECT 88.125 39.210 88.295 39.380 ;
        RECT 88.485 39.210 88.655 39.380 ;
        RECT 88.845 39.210 89.015 39.380 ;
        RECT 89.890 39.320 90.060 39.490 ;
        RECT 69.190 38.960 69.360 39.130 ;
        RECT 89.890 38.960 90.060 39.130 ;
        RECT 69.540 38.660 69.710 38.830 ;
        RECT 69.900 38.660 70.070 38.830 ;
        RECT 70.260 38.660 70.430 38.830 ;
        RECT 70.620 38.660 70.790 38.830 ;
        RECT 70.980 38.660 71.150 38.830 ;
        RECT 71.340 38.660 71.510 38.830 ;
        RECT 71.700 38.660 71.870 38.830 ;
        RECT 72.060 38.660 72.230 38.830 ;
        RECT 72.420 38.660 72.590 38.830 ;
        RECT 72.780 38.660 72.950 38.830 ;
        RECT 73.140 38.660 73.310 38.830 ;
        RECT 73.500 38.660 73.670 38.830 ;
        RECT 73.860 38.660 74.030 38.830 ;
        RECT 74.220 38.660 74.390 38.830 ;
        RECT 74.580 38.660 74.750 38.830 ;
        RECT 74.940 38.660 75.110 38.830 ;
        RECT 75.300 38.660 75.470 38.830 ;
        RECT 75.660 38.660 75.830 38.830 ;
        RECT 76.020 38.660 76.190 38.830 ;
        RECT 76.380 38.660 76.550 38.830 ;
        RECT 76.740 38.660 76.910 38.830 ;
        RECT 77.100 38.660 77.270 38.830 ;
        RECT 77.460 38.660 77.630 38.830 ;
        RECT 77.820 38.660 77.990 38.830 ;
        RECT 78.180 38.660 78.350 38.830 ;
        RECT 78.540 38.660 78.710 38.830 ;
        RECT 78.900 38.660 79.070 38.830 ;
        RECT 79.260 38.660 79.430 38.830 ;
        RECT 79.620 38.660 79.790 38.830 ;
        RECT 79.980 38.660 80.150 38.830 ;
        RECT 80.340 38.660 80.510 38.830 ;
        RECT 80.700 38.660 80.870 38.830 ;
        RECT 81.060 38.660 81.230 38.830 ;
        RECT 81.420 38.660 81.590 38.830 ;
        RECT 81.780 38.660 81.950 38.830 ;
        RECT 82.140 38.660 82.310 38.830 ;
        RECT 82.500 38.660 82.670 38.830 ;
        RECT 82.860 38.660 83.030 38.830 ;
        RECT 83.220 38.660 83.390 38.830 ;
        RECT 83.580 38.660 83.750 38.830 ;
        RECT 83.940 38.660 84.110 38.830 ;
        RECT 84.300 38.660 84.470 38.830 ;
        RECT 84.660 38.660 84.830 38.830 ;
        RECT 85.020 38.660 85.190 38.830 ;
        RECT 85.380 38.660 85.550 38.830 ;
        RECT 85.740 38.660 85.910 38.830 ;
        RECT 86.100 38.660 86.270 38.830 ;
        RECT 86.460 38.660 86.630 38.830 ;
        RECT 86.820 38.660 86.990 38.830 ;
        RECT 87.180 38.660 87.350 38.830 ;
        RECT 87.540 38.660 87.710 38.830 ;
        RECT 87.900 38.660 88.070 38.830 ;
        RECT 88.260 38.660 88.430 38.830 ;
        RECT 88.620 38.660 88.790 38.830 ;
        RECT 88.980 38.660 89.150 38.830 ;
        RECT 89.340 38.660 89.510 38.830 ;
        RECT 125.160 37.915 125.330 38.085 ;
        RECT 125.520 37.915 125.690 38.085 ;
        RECT 125.880 37.915 126.050 38.085 ;
        RECT 126.240 37.915 126.410 38.085 ;
        RECT 126.600 37.915 126.770 38.085 ;
        RECT 126.960 37.915 127.130 38.085 ;
        RECT 127.320 37.915 127.490 38.085 ;
        RECT 127.680 37.915 127.850 38.085 ;
        RECT 128.040 37.915 128.210 38.085 ;
        RECT 128.400 37.915 128.570 38.085 ;
        RECT 128.760 37.915 128.930 38.085 ;
        RECT 129.120 37.915 129.290 38.085 ;
        RECT 124.810 37.615 124.980 37.785 ;
        RECT 129.590 37.615 129.760 37.785 ;
        RECT 124.810 37.255 124.980 37.425 ;
        RECT 125.730 37.365 125.900 37.535 ;
        RECT 126.090 37.365 126.260 37.535 ;
        RECT 126.590 37.365 126.760 37.535 ;
        RECT 126.950 37.365 127.120 37.535 ;
        RECT 127.450 37.365 127.620 37.535 ;
        RECT 127.810 37.365 127.980 37.535 ;
        RECT 128.310 37.365 128.480 37.535 ;
        RECT 128.670 37.365 128.840 37.535 ;
        RECT 65.050 37.030 65.220 37.200 ;
        RECT 65.410 37.030 65.580 37.200 ;
        RECT 65.770 37.030 65.940 37.200 ;
        RECT 66.130 37.030 66.300 37.200 ;
        RECT 66.490 37.030 66.660 37.200 ;
        RECT 66.850 37.030 67.020 37.200 ;
        RECT 67.210 37.030 67.380 37.200 ;
        RECT 67.570 37.030 67.740 37.200 ;
        RECT 67.930 37.030 68.100 37.200 ;
        RECT 68.290 37.030 68.460 37.200 ;
        RECT 68.650 37.030 68.820 37.200 ;
        RECT 69.010 37.030 69.180 37.200 ;
        RECT 69.370 37.030 69.540 37.200 ;
        RECT 69.730 37.030 69.900 37.200 ;
        RECT 70.090 37.030 70.260 37.200 ;
        RECT 70.450 37.030 70.620 37.200 ;
        RECT 70.810 37.030 70.980 37.200 ;
        RECT 71.170 37.030 71.340 37.200 ;
        RECT 71.530 37.030 71.700 37.200 ;
        RECT 71.890 37.030 72.060 37.200 ;
        RECT 72.250 37.030 72.420 37.200 ;
        RECT 72.610 37.030 72.780 37.200 ;
        RECT 72.970 37.030 73.140 37.200 ;
        RECT 73.330 37.030 73.500 37.200 ;
        RECT 73.690 37.030 73.860 37.200 ;
        RECT 74.050 37.030 74.220 37.200 ;
        RECT 74.410 37.030 74.580 37.200 ;
        RECT 74.770 37.030 74.940 37.200 ;
        RECT 75.130 37.030 75.300 37.200 ;
        RECT 75.490 37.030 75.660 37.200 ;
        RECT 75.850 37.030 76.020 37.200 ;
        RECT 76.210 37.030 76.380 37.200 ;
        RECT 76.570 37.030 76.740 37.200 ;
        RECT 76.930 37.030 77.100 37.200 ;
        RECT 77.290 37.030 77.460 37.200 ;
        RECT 77.650 37.030 77.820 37.200 ;
        RECT 78.010 37.030 78.180 37.200 ;
        RECT 78.370 37.030 78.540 37.200 ;
        RECT 78.730 37.030 78.900 37.200 ;
        RECT 79.090 37.030 79.260 37.200 ;
        RECT 79.450 37.030 79.620 37.200 ;
        RECT 79.810 37.030 79.980 37.200 ;
        RECT 80.170 37.030 80.340 37.200 ;
        RECT 80.530 37.030 80.700 37.200 ;
        RECT 80.890 37.030 81.060 37.200 ;
        RECT 81.250 37.030 81.420 37.200 ;
        RECT 81.610 37.030 81.780 37.200 ;
        RECT 81.970 37.030 82.140 37.200 ;
        RECT 82.330 37.030 82.500 37.200 ;
        RECT 82.690 37.030 82.860 37.200 ;
        RECT 83.050 37.030 83.220 37.200 ;
        RECT 83.410 37.030 83.580 37.200 ;
        RECT 83.770 37.030 83.940 37.200 ;
        RECT 84.130 37.030 84.300 37.200 ;
        RECT 84.490 37.030 84.660 37.200 ;
        RECT 84.850 37.030 85.020 37.200 ;
        RECT 85.210 37.030 85.380 37.200 ;
        RECT 85.570 37.030 85.740 37.200 ;
        RECT 85.930 37.030 86.100 37.200 ;
        RECT 86.290 37.030 86.460 37.200 ;
        RECT 86.650 37.030 86.820 37.200 ;
        RECT 87.010 37.030 87.180 37.200 ;
        RECT 87.370 37.030 87.540 37.200 ;
        RECT 87.730 37.030 87.900 37.200 ;
        RECT 88.090 37.030 88.260 37.200 ;
        RECT 88.450 37.030 88.620 37.200 ;
        RECT 88.810 37.030 88.980 37.200 ;
        RECT 89.170 37.030 89.340 37.200 ;
        RECT 89.530 37.030 89.700 37.200 ;
        RECT 89.890 37.030 90.060 37.200 ;
        RECT 90.250 37.030 90.420 37.200 ;
        RECT 90.610 37.030 90.780 37.200 ;
        RECT 90.970 37.030 91.140 37.200 ;
        RECT 91.330 37.030 91.500 37.200 ;
        RECT 91.690 37.030 91.860 37.200 ;
        RECT 92.050 37.030 92.220 37.200 ;
        RECT 92.410 37.030 92.580 37.200 ;
        RECT 92.770 37.030 92.940 37.200 ;
        RECT 93.130 37.030 93.300 37.200 ;
        RECT 93.490 37.030 93.660 37.200 ;
        RECT 93.850 37.030 94.020 37.200 ;
        RECT 64.700 36.640 64.870 36.810 ;
        RECT 64.700 36.280 64.870 36.450 ;
        RECT 68.310 36.480 68.480 36.650 ;
        RECT 68.670 36.480 68.840 36.650 ;
        RECT 69.030 36.480 69.200 36.650 ;
        RECT 69.390 36.480 69.560 36.650 ;
        RECT 69.750 36.480 69.920 36.650 ;
        RECT 70.590 36.480 70.760 36.650 ;
        RECT 70.950 36.480 71.120 36.650 ;
        RECT 71.310 36.480 71.480 36.650 ;
        RECT 71.670 36.480 71.840 36.650 ;
        RECT 72.030 36.480 72.200 36.650 ;
        RECT 72.870 36.480 73.040 36.650 ;
        RECT 73.230 36.480 73.400 36.650 ;
        RECT 73.590 36.480 73.760 36.650 ;
        RECT 73.950 36.480 74.120 36.650 ;
        RECT 74.310 36.480 74.480 36.650 ;
        RECT 75.150 36.480 75.320 36.650 ;
        RECT 75.510 36.480 75.680 36.650 ;
        RECT 75.870 36.480 76.040 36.650 ;
        RECT 76.230 36.480 76.400 36.650 ;
        RECT 76.590 36.480 76.760 36.650 ;
        RECT 77.395 36.480 77.565 36.650 ;
        RECT 77.755 36.480 77.925 36.650 ;
        RECT 78.115 36.480 78.285 36.650 ;
        RECT 78.475 36.480 78.645 36.650 ;
        RECT 78.835 36.480 79.005 36.650 ;
        RECT 79.195 36.480 79.365 36.650 ;
        RECT 79.955 36.480 80.125 36.650 ;
        RECT 80.315 36.480 80.485 36.650 ;
        RECT 80.675 36.480 80.845 36.650 ;
        RECT 81.035 36.480 81.205 36.650 ;
        RECT 81.395 36.480 81.565 36.650 ;
        RECT 81.755 36.480 81.925 36.650 ;
        RECT 82.550 36.480 82.720 36.650 ;
        RECT 82.910 36.480 83.080 36.650 ;
        RECT 83.270 36.480 83.440 36.650 ;
        RECT 83.630 36.480 83.800 36.650 ;
        RECT 83.990 36.480 84.160 36.650 ;
        RECT 84.830 36.480 85.000 36.650 ;
        RECT 85.190 36.480 85.360 36.650 ;
        RECT 85.550 36.480 85.720 36.650 ;
        RECT 85.910 36.480 86.080 36.650 ;
        RECT 86.270 36.480 86.440 36.650 ;
        RECT 87.110 36.480 87.280 36.650 ;
        RECT 87.470 36.480 87.640 36.650 ;
        RECT 87.830 36.480 88.000 36.650 ;
        RECT 88.190 36.480 88.360 36.650 ;
        RECT 88.550 36.480 88.720 36.650 ;
        RECT 89.390 36.480 89.560 36.650 ;
        RECT 89.750 36.480 89.920 36.650 ;
        RECT 90.110 36.480 90.280 36.650 ;
        RECT 90.470 36.480 90.640 36.650 ;
        RECT 90.830 36.480 91.000 36.650 ;
        RECT 94.440 36.640 94.610 36.810 ;
        RECT 94.440 36.280 94.610 36.450 ;
        RECT 64.700 35.920 64.870 36.090 ;
        RECT 65.330 35.895 65.500 36.065 ;
        RECT 66.610 35.895 66.780 36.065 ;
        RECT 67.890 35.895 68.060 36.065 ;
        RECT 70.170 35.895 70.340 36.065 ;
        RECT 72.450 35.895 72.620 36.065 ;
        RECT 74.730 35.895 74.900 36.065 ;
        RECT 77.010 35.895 77.180 36.065 ;
        RECT 78.290 35.895 78.460 36.065 ;
        RECT 79.570 35.895 79.740 36.065 ;
        RECT 80.850 35.895 81.020 36.065 ;
        RECT 82.130 35.895 82.300 36.065 ;
        RECT 84.410 35.895 84.580 36.065 ;
        RECT 86.690 35.895 86.860 36.065 ;
        RECT 88.970 35.895 89.140 36.065 ;
        RECT 91.250 35.895 91.420 36.065 ;
        RECT 92.530 35.895 92.700 36.065 ;
        RECT 93.810 35.895 93.980 36.065 ;
        RECT 94.440 35.920 94.610 36.090 ;
        RECT 64.700 35.560 64.870 35.730 ;
        RECT 94.440 35.560 94.610 35.730 ;
        RECT 64.700 35.200 64.870 35.370 ;
        RECT 65.715 35.310 65.885 35.480 ;
        RECT 66.075 35.310 66.245 35.480 ;
        RECT 66.435 35.310 66.605 35.480 ;
        RECT 66.795 35.310 66.965 35.480 ;
        RECT 67.155 35.310 67.325 35.480 ;
        RECT 67.515 35.310 67.685 35.480 ;
        RECT 68.310 35.310 68.480 35.480 ;
        RECT 68.670 35.310 68.840 35.480 ;
        RECT 69.030 35.310 69.200 35.480 ;
        RECT 69.390 35.310 69.560 35.480 ;
        RECT 69.750 35.310 69.920 35.480 ;
        RECT 70.590 35.310 70.760 35.480 ;
        RECT 70.950 35.310 71.120 35.480 ;
        RECT 71.310 35.310 71.480 35.480 ;
        RECT 71.670 35.310 71.840 35.480 ;
        RECT 72.030 35.310 72.200 35.480 ;
        RECT 72.870 35.310 73.040 35.480 ;
        RECT 73.230 35.310 73.400 35.480 ;
        RECT 73.590 35.310 73.760 35.480 ;
        RECT 73.950 35.310 74.120 35.480 ;
        RECT 74.310 35.310 74.480 35.480 ;
        RECT 75.150 35.310 75.320 35.480 ;
        RECT 75.510 35.310 75.680 35.480 ;
        RECT 75.870 35.310 76.040 35.480 ;
        RECT 76.230 35.310 76.400 35.480 ;
        RECT 76.590 35.310 76.760 35.480 ;
        RECT 77.395 35.310 77.565 35.480 ;
        RECT 77.755 35.310 77.925 35.480 ;
        RECT 78.115 35.310 78.285 35.480 ;
        RECT 78.475 35.310 78.645 35.480 ;
        RECT 78.835 35.310 79.005 35.480 ;
        RECT 79.195 35.310 79.365 35.480 ;
        RECT 79.955 35.310 80.125 35.480 ;
        RECT 80.315 35.310 80.485 35.480 ;
        RECT 80.675 35.310 80.845 35.480 ;
        RECT 81.035 35.310 81.205 35.480 ;
        RECT 81.395 35.310 81.565 35.480 ;
        RECT 81.755 35.310 81.925 35.480 ;
        RECT 82.550 35.310 82.720 35.480 ;
        RECT 82.910 35.310 83.080 35.480 ;
        RECT 83.270 35.310 83.440 35.480 ;
        RECT 83.630 35.310 83.800 35.480 ;
        RECT 83.990 35.310 84.160 35.480 ;
        RECT 84.830 35.310 85.000 35.480 ;
        RECT 85.190 35.310 85.360 35.480 ;
        RECT 85.550 35.310 85.720 35.480 ;
        RECT 85.910 35.310 86.080 35.480 ;
        RECT 86.270 35.310 86.440 35.480 ;
        RECT 87.110 35.310 87.280 35.480 ;
        RECT 87.470 35.310 87.640 35.480 ;
        RECT 87.830 35.310 88.000 35.480 ;
        RECT 88.190 35.310 88.360 35.480 ;
        RECT 88.550 35.310 88.720 35.480 ;
        RECT 89.390 35.310 89.560 35.480 ;
        RECT 89.750 35.310 89.920 35.480 ;
        RECT 90.110 35.310 90.280 35.480 ;
        RECT 90.470 35.310 90.640 35.480 ;
        RECT 90.830 35.310 91.000 35.480 ;
        RECT 91.635 35.310 91.805 35.480 ;
        RECT 91.995 35.310 92.165 35.480 ;
        RECT 92.355 35.310 92.525 35.480 ;
        RECT 92.715 35.310 92.885 35.480 ;
        RECT 93.075 35.310 93.245 35.480 ;
        RECT 93.435 35.310 93.605 35.480 ;
        RECT 64.700 34.840 64.870 35.010 ;
        RECT 64.700 34.480 64.870 34.650 ;
        RECT 64.700 34.120 64.870 34.290 ;
        RECT 94.440 35.200 94.610 35.370 ;
        RECT 129.590 37.255 129.760 37.425 ;
        RECT 124.810 36.895 124.980 37.065 ;
        RECT 124.810 36.535 124.980 36.705 ;
        RECT 124.810 36.175 124.980 36.345 ;
        RECT 125.480 36.710 125.650 36.880 ;
        RECT 125.480 36.350 125.650 36.520 ;
        RECT 125.910 36.710 126.080 36.880 ;
        RECT 125.910 36.350 126.080 36.520 ;
        RECT 126.340 36.710 126.510 36.880 ;
        RECT 126.340 36.350 126.510 36.520 ;
        RECT 126.770 36.710 126.940 36.880 ;
        RECT 126.770 36.350 126.940 36.520 ;
        RECT 127.200 36.710 127.370 36.880 ;
        RECT 127.200 36.350 127.370 36.520 ;
        RECT 127.630 36.710 127.800 36.880 ;
        RECT 127.630 36.350 127.800 36.520 ;
        RECT 128.060 36.710 128.230 36.880 ;
        RECT 128.060 36.350 128.230 36.520 ;
        RECT 128.490 36.710 128.660 36.880 ;
        RECT 128.490 36.350 128.660 36.520 ;
        RECT 128.920 36.710 129.090 36.880 ;
        RECT 128.920 36.350 129.090 36.520 ;
        RECT 129.590 36.895 129.760 37.065 ;
        RECT 129.590 36.535 129.760 36.705 ;
        RECT 129.590 36.175 129.760 36.345 ;
        RECT 124.810 35.815 124.980 35.985 ;
        RECT 125.730 35.695 125.900 35.865 ;
        RECT 126.090 35.695 126.260 35.865 ;
        RECT 126.590 35.695 126.760 35.865 ;
        RECT 126.950 35.695 127.120 35.865 ;
        RECT 127.450 35.695 127.620 35.865 ;
        RECT 127.810 35.695 127.980 35.865 ;
        RECT 128.310 35.695 128.480 35.865 ;
        RECT 128.670 35.695 128.840 35.865 ;
        RECT 129.590 35.815 129.760 35.985 ;
        RECT 135.470 37.575 135.640 37.745 ;
        RECT 135.830 37.575 136.000 37.745 ;
        RECT 136.190 37.575 136.360 37.745 ;
        RECT 136.550 37.575 136.720 37.745 ;
        RECT 136.910 37.575 137.080 37.745 ;
        RECT 137.270 37.575 137.440 37.745 ;
        RECT 137.630 37.575 137.800 37.745 ;
        RECT 137.990 37.575 138.160 37.745 ;
        RECT 138.350 37.575 138.520 37.745 ;
        RECT 138.710 37.575 138.880 37.745 ;
        RECT 139.070 37.575 139.240 37.745 ;
        RECT 139.430 37.575 139.600 37.745 ;
        RECT 139.790 37.575 139.960 37.745 ;
        RECT 140.150 37.575 140.320 37.745 ;
        RECT 140.510 37.575 140.680 37.745 ;
        RECT 140.870 37.575 141.040 37.745 ;
        RECT 141.230 37.575 141.400 37.745 ;
        RECT 141.590 37.575 141.760 37.745 ;
        RECT 141.950 37.575 142.120 37.745 ;
        RECT 142.310 37.575 142.480 37.745 ;
        RECT 142.670 37.575 142.840 37.745 ;
        RECT 143.030 37.575 143.200 37.745 ;
        RECT 143.390 37.575 143.560 37.745 ;
        RECT 143.750 37.575 143.920 37.745 ;
        RECT 135.120 37.275 135.290 37.445 ;
        RECT 144.200 37.275 144.370 37.445 ;
        RECT 135.120 36.915 135.290 37.085 ;
        RECT 135.120 36.555 135.290 36.725 ;
        RECT 135.120 36.195 135.290 36.365 ;
        RECT 135.790 36.735 135.960 36.905 ;
        RECT 135.790 36.375 135.960 36.545 ;
        RECT 136.220 36.735 136.390 36.905 ;
        RECT 136.220 36.375 136.390 36.545 ;
        RECT 136.650 36.735 136.820 36.905 ;
        RECT 136.650 36.375 136.820 36.545 ;
        RECT 137.080 36.735 137.250 36.905 ;
        RECT 137.080 36.375 137.250 36.545 ;
        RECT 137.510 36.735 137.680 36.905 ;
        RECT 137.510 36.375 137.680 36.545 ;
        RECT 137.940 36.735 138.110 36.905 ;
        RECT 137.940 36.375 138.110 36.545 ;
        RECT 138.370 36.735 138.540 36.905 ;
        RECT 138.370 36.375 138.540 36.545 ;
        RECT 138.800 36.735 138.970 36.905 ;
        RECT 138.800 36.375 138.970 36.545 ;
        RECT 139.230 36.735 139.400 36.905 ;
        RECT 139.230 36.375 139.400 36.545 ;
        RECT 139.660 36.735 139.830 36.905 ;
        RECT 139.660 36.375 139.830 36.545 ;
        RECT 140.090 36.735 140.260 36.905 ;
        RECT 140.090 36.375 140.260 36.545 ;
        RECT 140.520 36.735 140.690 36.905 ;
        RECT 140.520 36.375 140.690 36.545 ;
        RECT 140.950 36.735 141.120 36.905 ;
        RECT 140.950 36.375 141.120 36.545 ;
        RECT 141.380 36.735 141.550 36.905 ;
        RECT 141.380 36.375 141.550 36.545 ;
        RECT 141.810 36.735 141.980 36.905 ;
        RECT 141.810 36.375 141.980 36.545 ;
        RECT 142.240 36.735 142.410 36.905 ;
        RECT 142.240 36.375 142.410 36.545 ;
        RECT 142.670 36.735 142.840 36.905 ;
        RECT 142.670 36.375 142.840 36.545 ;
        RECT 143.100 36.735 143.270 36.905 ;
        RECT 143.100 36.375 143.270 36.545 ;
        RECT 143.530 36.735 143.700 36.905 ;
        RECT 143.530 36.375 143.700 36.545 ;
        RECT 144.200 36.915 144.370 37.085 ;
        RECT 144.200 36.555 144.370 36.725 ;
        RECT 144.200 36.195 144.370 36.365 ;
        RECT 135.120 35.835 135.290 36.005 ;
        RECT 135.120 35.475 135.290 35.645 ;
        RECT 136.040 35.720 136.210 35.890 ;
        RECT 136.400 35.720 136.570 35.890 ;
        RECT 136.900 35.720 137.070 35.890 ;
        RECT 137.260 35.720 137.430 35.890 ;
        RECT 137.760 35.720 137.930 35.890 ;
        RECT 138.120 35.720 138.290 35.890 ;
        RECT 138.620 35.720 138.790 35.890 ;
        RECT 138.980 35.720 139.150 35.890 ;
        RECT 139.480 35.720 139.650 35.890 ;
        RECT 139.840 35.720 140.010 35.890 ;
        RECT 140.340 35.720 140.510 35.890 ;
        RECT 140.700 35.720 140.870 35.890 ;
        RECT 141.200 35.720 141.370 35.890 ;
        RECT 141.560 35.720 141.730 35.890 ;
        RECT 142.060 35.720 142.230 35.890 ;
        RECT 142.420 35.720 142.590 35.890 ;
        RECT 142.920 35.720 143.090 35.890 ;
        RECT 143.280 35.720 143.450 35.890 ;
        RECT 144.200 35.835 144.370 36.005 ;
        RECT 144.200 35.475 144.370 35.645 ;
        RECT 94.440 34.840 94.610 35.010 ;
        RECT 94.440 34.480 94.610 34.650 ;
        RECT 94.440 34.120 94.610 34.290 ;
        RECT 64.700 33.760 64.870 33.930 ;
        RECT 66.115 33.740 66.285 33.910 ;
        RECT 66.475 33.740 66.645 33.910 ;
        RECT 66.835 33.740 67.005 33.910 ;
        RECT 67.195 33.740 67.365 33.910 ;
        RECT 67.555 33.740 67.725 33.910 ;
        RECT 67.915 33.740 68.085 33.910 ;
        RECT 68.275 33.740 68.445 33.910 ;
        RECT 68.635 33.740 68.805 33.910 ;
        RECT 69.395 33.740 69.565 33.910 ;
        RECT 69.755 33.740 69.925 33.910 ;
        RECT 70.115 33.740 70.285 33.910 ;
        RECT 70.475 33.740 70.645 33.910 ;
        RECT 70.835 33.740 71.005 33.910 ;
        RECT 71.195 33.740 71.365 33.910 ;
        RECT 71.555 33.740 71.725 33.910 ;
        RECT 71.915 33.740 72.085 33.910 ;
        RECT 87.235 33.740 87.405 33.910 ;
        RECT 87.595 33.740 87.765 33.910 ;
        RECT 87.955 33.740 88.125 33.910 ;
        RECT 88.315 33.740 88.485 33.910 ;
        RECT 88.675 33.740 88.845 33.910 ;
        RECT 89.035 33.740 89.205 33.910 ;
        RECT 89.395 33.740 89.565 33.910 ;
        RECT 89.755 33.740 89.925 33.910 ;
        RECT 90.515 33.740 90.685 33.910 ;
        RECT 90.875 33.740 91.045 33.910 ;
        RECT 91.235 33.740 91.405 33.910 ;
        RECT 91.595 33.740 91.765 33.910 ;
        RECT 91.955 33.740 92.125 33.910 ;
        RECT 92.315 33.740 92.485 33.910 ;
        RECT 92.675 33.740 92.845 33.910 ;
        RECT 93.035 33.740 93.205 33.910 ;
        RECT 94.440 33.760 94.610 33.930 ;
        RECT 64.700 33.400 64.870 33.570 ;
        RECT 64.700 33.040 64.870 33.210 ;
        RECT 65.730 33.155 65.900 33.325 ;
        RECT 69.010 33.155 69.180 33.325 ;
        RECT 72.290 33.155 72.460 33.325 ;
        RECT 79.570 33.155 79.740 33.325 ;
        RECT 86.850 33.155 87.020 33.325 ;
        RECT 90.130 33.155 90.300 33.325 ;
        RECT 93.410 33.155 93.580 33.325 ;
        RECT 94.440 33.400 94.610 33.570 ;
        RECT 94.440 33.040 94.610 33.210 ;
        RECT 64.700 32.680 64.870 32.850 ;
        RECT 66.115 32.570 66.285 32.740 ;
        RECT 66.475 32.570 66.645 32.740 ;
        RECT 66.835 32.570 67.005 32.740 ;
        RECT 67.195 32.570 67.365 32.740 ;
        RECT 67.555 32.570 67.725 32.740 ;
        RECT 67.915 32.570 68.085 32.740 ;
        RECT 68.275 32.570 68.445 32.740 ;
        RECT 68.635 32.570 68.805 32.740 ;
        RECT 69.395 32.570 69.565 32.740 ;
        RECT 69.755 32.570 69.925 32.740 ;
        RECT 70.115 32.570 70.285 32.740 ;
        RECT 70.475 32.570 70.645 32.740 ;
        RECT 70.835 32.570 71.005 32.740 ;
        RECT 71.195 32.570 71.365 32.740 ;
        RECT 71.555 32.570 71.725 32.740 ;
        RECT 71.915 32.570 72.085 32.740 ;
        RECT 72.690 32.570 72.860 32.740 ;
        RECT 73.050 32.570 73.220 32.740 ;
        RECT 73.410 32.570 73.580 32.740 ;
        RECT 73.770 32.570 73.940 32.740 ;
        RECT 74.130 32.570 74.300 32.740 ;
        RECT 74.490 32.570 74.660 32.740 ;
        RECT 74.850 32.570 75.020 32.740 ;
        RECT 75.210 32.570 75.380 32.740 ;
        RECT 75.570 32.570 75.740 32.740 ;
        RECT 75.930 32.570 76.100 32.740 ;
        RECT 76.290 32.570 76.460 32.740 ;
        RECT 76.650 32.570 76.820 32.740 ;
        RECT 77.010 32.570 77.180 32.740 ;
        RECT 77.370 32.570 77.540 32.740 ;
        RECT 77.730 32.570 77.900 32.740 ;
        RECT 78.090 32.570 78.260 32.740 ;
        RECT 78.450 32.570 78.620 32.740 ;
        RECT 78.810 32.570 78.980 32.740 ;
        RECT 79.170 32.570 79.340 32.740 ;
        RECT 79.970 32.570 80.140 32.740 ;
        RECT 80.330 32.570 80.500 32.740 ;
        RECT 80.690 32.570 80.860 32.740 ;
        RECT 81.050 32.570 81.220 32.740 ;
        RECT 81.410 32.570 81.580 32.740 ;
        RECT 81.770 32.570 81.940 32.740 ;
        RECT 82.130 32.570 82.300 32.740 ;
        RECT 82.490 32.570 82.660 32.740 ;
        RECT 82.850 32.570 83.020 32.740 ;
        RECT 83.210 32.570 83.380 32.740 ;
        RECT 83.570 32.570 83.740 32.740 ;
        RECT 83.930 32.570 84.100 32.740 ;
        RECT 84.290 32.570 84.460 32.740 ;
        RECT 84.650 32.570 84.820 32.740 ;
        RECT 85.010 32.570 85.180 32.740 ;
        RECT 85.370 32.570 85.540 32.740 ;
        RECT 85.730 32.570 85.900 32.740 ;
        RECT 86.090 32.570 86.260 32.740 ;
        RECT 86.450 32.570 86.620 32.740 ;
        RECT 87.235 32.570 87.405 32.740 ;
        RECT 87.595 32.570 87.765 32.740 ;
        RECT 87.955 32.570 88.125 32.740 ;
        RECT 88.315 32.570 88.485 32.740 ;
        RECT 88.675 32.570 88.845 32.740 ;
        RECT 89.035 32.570 89.205 32.740 ;
        RECT 89.395 32.570 89.565 32.740 ;
        RECT 89.755 32.570 89.925 32.740 ;
        RECT 90.515 32.570 90.685 32.740 ;
        RECT 90.875 32.570 91.045 32.740 ;
        RECT 91.235 32.570 91.405 32.740 ;
        RECT 91.595 32.570 91.765 32.740 ;
        RECT 91.955 32.570 92.125 32.740 ;
        RECT 92.315 32.570 92.485 32.740 ;
        RECT 92.675 32.570 92.845 32.740 ;
        RECT 93.035 32.570 93.205 32.740 ;
        RECT 94.440 32.680 94.610 32.850 ;
        RECT 64.700 32.320 64.870 32.490 ;
        RECT 94.440 32.320 94.610 32.490 ;
        RECT 65.050 32.020 65.220 32.190 ;
        RECT 65.410 32.020 65.580 32.190 ;
        RECT 65.770 32.020 65.940 32.190 ;
        RECT 66.130 32.020 66.300 32.190 ;
        RECT 66.490 32.020 66.660 32.190 ;
        RECT 66.850 32.020 67.020 32.190 ;
        RECT 67.210 32.020 67.380 32.190 ;
        RECT 67.570 32.020 67.740 32.190 ;
        RECT 67.930 32.020 68.100 32.190 ;
        RECT 68.290 32.020 68.460 32.190 ;
        RECT 68.650 32.020 68.820 32.190 ;
        RECT 69.010 32.020 69.180 32.190 ;
        RECT 69.370 32.020 69.540 32.190 ;
        RECT 69.730 32.020 69.900 32.190 ;
        RECT 70.090 32.020 70.260 32.190 ;
        RECT 70.450 32.020 70.620 32.190 ;
        RECT 70.810 32.020 70.980 32.190 ;
        RECT 71.170 32.020 71.340 32.190 ;
        RECT 71.530 32.020 71.700 32.190 ;
        RECT 71.890 32.020 72.060 32.190 ;
        RECT 72.250 32.020 72.420 32.190 ;
        RECT 72.610 32.020 72.780 32.190 ;
        RECT 72.970 32.020 73.140 32.190 ;
        RECT 73.330 32.020 73.500 32.190 ;
        RECT 73.690 32.020 73.860 32.190 ;
        RECT 74.050 32.020 74.220 32.190 ;
        RECT 74.410 32.020 74.580 32.190 ;
        RECT 74.770 32.020 74.940 32.190 ;
        RECT 75.130 32.020 75.300 32.190 ;
        RECT 75.490 32.020 75.660 32.190 ;
        RECT 75.850 32.020 76.020 32.190 ;
        RECT 76.210 32.020 76.380 32.190 ;
        RECT 76.570 32.020 76.740 32.190 ;
        RECT 76.930 32.020 77.100 32.190 ;
        RECT 77.290 32.020 77.460 32.190 ;
        RECT 77.650 32.020 77.820 32.190 ;
        RECT 78.010 32.020 78.180 32.190 ;
        RECT 78.370 32.020 78.540 32.190 ;
        RECT 78.730 32.020 78.900 32.190 ;
        RECT 79.090 32.020 79.260 32.190 ;
        RECT 79.450 32.020 79.620 32.190 ;
        RECT 79.810 32.020 79.980 32.190 ;
        RECT 80.170 32.020 80.340 32.190 ;
        RECT 80.530 32.020 80.700 32.190 ;
        RECT 80.890 32.020 81.060 32.190 ;
        RECT 81.250 32.020 81.420 32.190 ;
        RECT 81.610 32.020 81.780 32.190 ;
        RECT 81.970 32.020 82.140 32.190 ;
        RECT 82.330 32.020 82.500 32.190 ;
        RECT 82.690 32.020 82.860 32.190 ;
        RECT 83.050 32.020 83.220 32.190 ;
        RECT 83.410 32.020 83.580 32.190 ;
        RECT 83.770 32.020 83.940 32.190 ;
        RECT 84.130 32.020 84.300 32.190 ;
        RECT 84.490 32.020 84.660 32.190 ;
        RECT 84.850 32.020 85.020 32.190 ;
        RECT 85.210 32.020 85.380 32.190 ;
        RECT 85.570 32.020 85.740 32.190 ;
        RECT 85.930 32.020 86.100 32.190 ;
        RECT 86.290 32.020 86.460 32.190 ;
        RECT 86.650 32.020 86.820 32.190 ;
        RECT 87.010 32.020 87.180 32.190 ;
        RECT 87.370 32.020 87.540 32.190 ;
        RECT 87.730 32.020 87.900 32.190 ;
        RECT 88.090 32.020 88.260 32.190 ;
        RECT 88.450 32.020 88.620 32.190 ;
        RECT 88.810 32.020 88.980 32.190 ;
        RECT 89.170 32.020 89.340 32.190 ;
        RECT 89.530 32.020 89.700 32.190 ;
        RECT 89.890 32.020 90.060 32.190 ;
        RECT 90.250 32.020 90.420 32.190 ;
        RECT 90.610 32.020 90.780 32.190 ;
        RECT 90.970 32.020 91.140 32.190 ;
        RECT 91.330 32.020 91.500 32.190 ;
        RECT 91.690 32.020 91.860 32.190 ;
        RECT 92.050 32.020 92.220 32.190 ;
        RECT 92.410 32.020 92.580 32.190 ;
        RECT 92.770 32.020 92.940 32.190 ;
        RECT 93.130 32.020 93.300 32.190 ;
        RECT 93.490 32.020 93.660 32.190 ;
        RECT 93.850 32.020 94.020 32.190 ;
        RECT 124.810 34.095 124.980 34.265 ;
        RECT 125.730 34.065 125.900 34.235 ;
        RECT 126.090 34.065 126.260 34.235 ;
        RECT 126.590 34.065 126.760 34.235 ;
        RECT 126.950 34.065 127.120 34.235 ;
        RECT 127.450 34.065 127.620 34.235 ;
        RECT 127.810 34.065 127.980 34.235 ;
        RECT 128.310 34.065 128.480 34.235 ;
        RECT 128.670 34.065 128.840 34.235 ;
        RECT 129.590 34.095 129.760 34.265 ;
        RECT 124.810 33.735 124.980 33.905 ;
        RECT 124.810 33.375 124.980 33.545 ;
        RECT 124.810 33.015 124.980 33.185 ;
        RECT 124.810 32.655 124.980 32.825 ;
        RECT 125.480 33.410 125.650 33.580 ;
        RECT 125.480 33.050 125.650 33.220 ;
        RECT 125.910 33.410 126.080 33.580 ;
        RECT 125.910 33.050 126.080 33.220 ;
        RECT 126.340 33.410 126.510 33.580 ;
        RECT 126.340 33.050 126.510 33.220 ;
        RECT 126.770 33.410 126.940 33.580 ;
        RECT 126.770 33.050 126.940 33.220 ;
        RECT 127.200 33.410 127.370 33.580 ;
        RECT 127.200 33.050 127.370 33.220 ;
        RECT 127.630 33.410 127.800 33.580 ;
        RECT 127.630 33.050 127.800 33.220 ;
        RECT 128.060 33.410 128.230 33.580 ;
        RECT 128.060 33.050 128.230 33.220 ;
        RECT 128.490 33.410 128.660 33.580 ;
        RECT 128.490 33.050 128.660 33.220 ;
        RECT 128.920 33.410 129.090 33.580 ;
        RECT 128.920 33.050 129.090 33.220 ;
        RECT 129.590 33.735 129.760 33.905 ;
        RECT 129.590 33.375 129.760 33.545 ;
        RECT 129.590 33.015 129.760 33.185 ;
        RECT 124.810 32.295 124.980 32.465 ;
        RECT 129.590 32.655 129.760 32.825 ;
        RECT 129.590 32.295 129.760 32.465 ;
        RECT 124.810 31.935 124.980 32.105 ;
        RECT 124.810 31.575 124.980 31.745 ;
        RECT 124.810 31.215 124.980 31.385 ;
        RECT 125.480 31.760 125.650 31.930 ;
        RECT 125.480 31.400 125.650 31.570 ;
        RECT 125.910 31.760 126.080 31.930 ;
        RECT 125.910 31.400 126.080 31.570 ;
        RECT 126.340 31.760 126.510 31.930 ;
        RECT 126.340 31.400 126.510 31.570 ;
        RECT 126.770 31.760 126.940 31.930 ;
        RECT 126.770 31.400 126.940 31.570 ;
        RECT 127.200 31.760 127.370 31.930 ;
        RECT 127.200 31.400 127.370 31.570 ;
        RECT 127.630 31.760 127.800 31.930 ;
        RECT 127.630 31.400 127.800 31.570 ;
        RECT 128.060 31.760 128.230 31.930 ;
        RECT 128.060 31.400 128.230 31.570 ;
        RECT 128.490 31.760 128.660 31.930 ;
        RECT 128.490 31.400 128.660 31.570 ;
        RECT 128.920 31.760 129.090 31.930 ;
        RECT 128.920 31.400 129.090 31.570 ;
        RECT 129.590 31.935 129.760 32.105 ;
        RECT 129.590 31.575 129.760 31.745 ;
        RECT 129.590 31.215 129.760 31.385 ;
        RECT 124.810 30.855 124.980 31.025 ;
        RECT 125.730 30.745 125.900 30.915 ;
        RECT 126.090 30.745 126.260 30.915 ;
        RECT 126.590 30.745 126.760 30.915 ;
        RECT 126.950 30.745 127.120 30.915 ;
        RECT 127.450 30.745 127.620 30.915 ;
        RECT 127.810 30.745 127.980 30.915 ;
        RECT 128.310 30.745 128.480 30.915 ;
        RECT 128.670 30.745 128.840 30.915 ;
        RECT 129.590 30.855 129.760 31.025 ;
        RECT 124.810 30.495 124.980 30.665 ;
        RECT 129.590 30.495 129.760 30.665 ;
        RECT 125.160 30.195 125.330 30.365 ;
        RECT 125.520 30.195 125.690 30.365 ;
        RECT 125.880 30.195 126.050 30.365 ;
        RECT 126.240 30.195 126.410 30.365 ;
        RECT 126.600 30.195 126.770 30.365 ;
        RECT 126.960 30.195 127.130 30.365 ;
        RECT 127.320 30.195 127.490 30.365 ;
        RECT 127.680 30.195 127.850 30.365 ;
        RECT 128.040 30.195 128.210 30.365 ;
        RECT 128.400 30.195 128.570 30.365 ;
        RECT 128.760 30.195 128.930 30.365 ;
        RECT 129.120 30.195 129.290 30.365 ;
        RECT 124.810 29.895 124.980 30.065 ;
        RECT 129.590 29.895 129.760 30.065 ;
        RECT 124.810 29.535 124.980 29.705 ;
        RECT 125.730 29.645 125.900 29.815 ;
        RECT 126.090 29.645 126.260 29.815 ;
        RECT 126.590 29.645 126.760 29.815 ;
        RECT 126.950 29.645 127.120 29.815 ;
        RECT 127.450 29.645 127.620 29.815 ;
        RECT 127.810 29.645 127.980 29.815 ;
        RECT 128.310 29.645 128.480 29.815 ;
        RECT 128.670 29.645 128.840 29.815 ;
        RECT 129.590 29.535 129.760 29.705 ;
        RECT 124.810 29.175 124.980 29.345 ;
        RECT 124.810 28.815 124.980 28.985 ;
        RECT 65.050 28.600 65.220 28.770 ;
        RECT 65.410 28.600 65.580 28.770 ;
        RECT 65.770 28.600 65.940 28.770 ;
        RECT 66.130 28.600 66.300 28.770 ;
        RECT 66.490 28.600 66.660 28.770 ;
        RECT 66.850 28.600 67.020 28.770 ;
        RECT 67.210 28.600 67.380 28.770 ;
        RECT 67.570 28.600 67.740 28.770 ;
        RECT 67.930 28.600 68.100 28.770 ;
        RECT 68.290 28.600 68.460 28.770 ;
        RECT 68.650 28.600 68.820 28.770 ;
        RECT 69.010 28.600 69.180 28.770 ;
        RECT 69.370 28.600 69.540 28.770 ;
        RECT 69.730 28.600 69.900 28.770 ;
        RECT 70.090 28.600 70.260 28.770 ;
        RECT 70.450 28.600 70.620 28.770 ;
        RECT 70.810 28.600 70.980 28.770 ;
        RECT 71.170 28.600 71.340 28.770 ;
        RECT 71.530 28.600 71.700 28.770 ;
        RECT 71.890 28.600 72.060 28.770 ;
        RECT 72.250 28.600 72.420 28.770 ;
        RECT 72.610 28.600 72.780 28.770 ;
        RECT 72.970 28.600 73.140 28.770 ;
        RECT 73.330 28.600 73.500 28.770 ;
        RECT 73.690 28.600 73.860 28.770 ;
        RECT 74.050 28.600 74.220 28.770 ;
        RECT 74.410 28.600 74.580 28.770 ;
        RECT 74.770 28.600 74.940 28.770 ;
        RECT 75.130 28.600 75.300 28.770 ;
        RECT 75.490 28.600 75.660 28.770 ;
        RECT 75.850 28.600 76.020 28.770 ;
        RECT 76.210 28.600 76.380 28.770 ;
        RECT 76.570 28.600 76.740 28.770 ;
        RECT 76.930 28.600 77.100 28.770 ;
        RECT 77.290 28.600 77.460 28.770 ;
        RECT 77.650 28.600 77.820 28.770 ;
        RECT 78.010 28.600 78.180 28.770 ;
        RECT 78.370 28.600 78.540 28.770 ;
        RECT 78.730 28.600 78.900 28.770 ;
        RECT 79.090 28.600 79.260 28.770 ;
        RECT 79.450 28.600 79.620 28.770 ;
        RECT 79.810 28.600 79.980 28.770 ;
        RECT 80.170 28.600 80.340 28.770 ;
        RECT 80.530 28.600 80.700 28.770 ;
        RECT 80.890 28.600 81.060 28.770 ;
        RECT 81.250 28.600 81.420 28.770 ;
        RECT 81.610 28.600 81.780 28.770 ;
        RECT 81.970 28.600 82.140 28.770 ;
        RECT 82.330 28.600 82.500 28.770 ;
        RECT 82.690 28.600 82.860 28.770 ;
        RECT 83.050 28.600 83.220 28.770 ;
        RECT 83.410 28.600 83.580 28.770 ;
        RECT 83.770 28.600 83.940 28.770 ;
        RECT 84.130 28.600 84.300 28.770 ;
        RECT 84.490 28.600 84.660 28.770 ;
        RECT 84.850 28.600 85.020 28.770 ;
        RECT 85.210 28.600 85.380 28.770 ;
        RECT 85.570 28.600 85.740 28.770 ;
        RECT 85.930 28.600 86.100 28.770 ;
        RECT 86.290 28.600 86.460 28.770 ;
        RECT 86.650 28.600 86.820 28.770 ;
        RECT 87.010 28.600 87.180 28.770 ;
        RECT 87.370 28.600 87.540 28.770 ;
        RECT 87.730 28.600 87.900 28.770 ;
        RECT 88.090 28.600 88.260 28.770 ;
        RECT 88.450 28.600 88.620 28.770 ;
        RECT 88.810 28.600 88.980 28.770 ;
        RECT 89.170 28.600 89.340 28.770 ;
        RECT 89.530 28.600 89.700 28.770 ;
        RECT 89.890 28.600 90.060 28.770 ;
        RECT 90.250 28.600 90.420 28.770 ;
        RECT 90.610 28.600 90.780 28.770 ;
        RECT 90.970 28.600 91.140 28.770 ;
        RECT 91.330 28.600 91.500 28.770 ;
        RECT 91.690 28.600 91.860 28.770 ;
        RECT 92.050 28.600 92.220 28.770 ;
        RECT 92.410 28.600 92.580 28.770 ;
        RECT 92.770 28.600 92.940 28.770 ;
        RECT 93.130 28.600 93.300 28.770 ;
        RECT 93.490 28.600 93.660 28.770 ;
        RECT 93.850 28.600 94.020 28.770 ;
        RECT 64.700 28.300 64.870 28.470 ;
        RECT 94.440 28.300 94.610 28.470 ;
        RECT 64.700 27.940 64.870 28.110 ;
        RECT 66.115 28.050 66.285 28.220 ;
        RECT 66.475 28.050 66.645 28.220 ;
        RECT 66.835 28.050 67.005 28.220 ;
        RECT 67.195 28.050 67.365 28.220 ;
        RECT 67.555 28.050 67.725 28.220 ;
        RECT 67.915 28.050 68.085 28.220 ;
        RECT 68.275 28.050 68.445 28.220 ;
        RECT 68.635 28.050 68.805 28.220 ;
        RECT 69.395 28.050 69.565 28.220 ;
        RECT 69.755 28.050 69.925 28.220 ;
        RECT 70.115 28.050 70.285 28.220 ;
        RECT 70.475 28.050 70.645 28.220 ;
        RECT 70.835 28.050 71.005 28.220 ;
        RECT 71.195 28.050 71.365 28.220 ;
        RECT 71.555 28.050 71.725 28.220 ;
        RECT 71.915 28.050 72.085 28.220 ;
        RECT 72.690 28.050 72.860 28.220 ;
        RECT 73.050 28.050 73.220 28.220 ;
        RECT 73.410 28.050 73.580 28.220 ;
        RECT 73.770 28.050 73.940 28.220 ;
        RECT 74.130 28.050 74.300 28.220 ;
        RECT 74.490 28.050 74.660 28.220 ;
        RECT 74.850 28.050 75.020 28.220 ;
        RECT 75.210 28.050 75.380 28.220 ;
        RECT 75.570 28.050 75.740 28.220 ;
        RECT 75.930 28.050 76.100 28.220 ;
        RECT 76.290 28.050 76.460 28.220 ;
        RECT 76.650 28.050 76.820 28.220 ;
        RECT 77.010 28.050 77.180 28.220 ;
        RECT 77.370 28.050 77.540 28.220 ;
        RECT 77.730 28.050 77.900 28.220 ;
        RECT 78.090 28.050 78.260 28.220 ;
        RECT 78.450 28.050 78.620 28.220 ;
        RECT 78.810 28.050 78.980 28.220 ;
        RECT 79.170 28.050 79.340 28.220 ;
        RECT 79.970 28.050 80.140 28.220 ;
        RECT 80.330 28.050 80.500 28.220 ;
        RECT 80.690 28.050 80.860 28.220 ;
        RECT 81.050 28.050 81.220 28.220 ;
        RECT 81.410 28.050 81.580 28.220 ;
        RECT 81.770 28.050 81.940 28.220 ;
        RECT 82.130 28.050 82.300 28.220 ;
        RECT 82.490 28.050 82.660 28.220 ;
        RECT 82.850 28.050 83.020 28.220 ;
        RECT 83.210 28.050 83.380 28.220 ;
        RECT 83.570 28.050 83.740 28.220 ;
        RECT 83.930 28.050 84.100 28.220 ;
        RECT 84.290 28.050 84.460 28.220 ;
        RECT 84.650 28.050 84.820 28.220 ;
        RECT 85.010 28.050 85.180 28.220 ;
        RECT 85.370 28.050 85.540 28.220 ;
        RECT 85.730 28.050 85.900 28.220 ;
        RECT 86.090 28.050 86.260 28.220 ;
        RECT 86.450 28.050 86.620 28.220 ;
        RECT 87.235 28.050 87.405 28.220 ;
        RECT 87.595 28.050 87.765 28.220 ;
        RECT 87.955 28.050 88.125 28.220 ;
        RECT 88.315 28.050 88.485 28.220 ;
        RECT 88.675 28.050 88.845 28.220 ;
        RECT 89.035 28.050 89.205 28.220 ;
        RECT 89.395 28.050 89.565 28.220 ;
        RECT 89.755 28.050 89.925 28.220 ;
        RECT 90.515 28.050 90.685 28.220 ;
        RECT 90.875 28.050 91.045 28.220 ;
        RECT 91.235 28.050 91.405 28.220 ;
        RECT 91.595 28.050 91.765 28.220 ;
        RECT 91.955 28.050 92.125 28.220 ;
        RECT 92.315 28.050 92.485 28.220 ;
        RECT 92.675 28.050 92.845 28.220 ;
        RECT 93.035 28.050 93.205 28.220 ;
        RECT 94.440 27.940 94.610 28.110 ;
        RECT 64.700 27.580 64.870 27.750 ;
        RECT 64.700 27.220 64.870 27.390 ;
        RECT 65.730 27.465 65.900 27.635 ;
        RECT 69.010 27.465 69.180 27.635 ;
        RECT 72.290 27.465 72.460 27.635 ;
        RECT 79.570 27.465 79.740 27.635 ;
        RECT 86.850 27.465 87.020 27.635 ;
        RECT 90.130 27.465 90.300 27.635 ;
        RECT 93.410 27.465 93.580 27.635 ;
        RECT 94.440 27.580 94.610 27.750 ;
        RECT 94.440 27.220 94.610 27.390 ;
        RECT 64.700 26.860 64.870 27.030 ;
        RECT 66.115 26.880 66.285 27.050 ;
        RECT 66.475 26.880 66.645 27.050 ;
        RECT 66.835 26.880 67.005 27.050 ;
        RECT 67.195 26.880 67.365 27.050 ;
        RECT 67.555 26.880 67.725 27.050 ;
        RECT 67.915 26.880 68.085 27.050 ;
        RECT 68.275 26.880 68.445 27.050 ;
        RECT 68.635 26.880 68.805 27.050 ;
        RECT 69.395 26.880 69.565 27.050 ;
        RECT 69.755 26.880 69.925 27.050 ;
        RECT 70.115 26.880 70.285 27.050 ;
        RECT 70.475 26.880 70.645 27.050 ;
        RECT 70.835 26.880 71.005 27.050 ;
        RECT 71.195 26.880 71.365 27.050 ;
        RECT 71.555 26.880 71.725 27.050 ;
        RECT 71.915 26.880 72.085 27.050 ;
        RECT 87.235 26.880 87.405 27.050 ;
        RECT 87.595 26.880 87.765 27.050 ;
        RECT 87.955 26.880 88.125 27.050 ;
        RECT 88.315 26.880 88.485 27.050 ;
        RECT 88.675 26.880 88.845 27.050 ;
        RECT 89.035 26.880 89.205 27.050 ;
        RECT 89.395 26.880 89.565 27.050 ;
        RECT 89.755 26.880 89.925 27.050 ;
        RECT 90.515 26.880 90.685 27.050 ;
        RECT 90.875 26.880 91.045 27.050 ;
        RECT 91.235 26.880 91.405 27.050 ;
        RECT 91.595 26.880 91.765 27.050 ;
        RECT 91.955 26.880 92.125 27.050 ;
        RECT 92.315 26.880 92.485 27.050 ;
        RECT 92.675 26.880 92.845 27.050 ;
        RECT 93.035 26.880 93.205 27.050 ;
        RECT 94.440 26.860 94.610 27.030 ;
        RECT 64.700 26.500 64.870 26.670 ;
        RECT 64.700 26.140 64.870 26.310 ;
        RECT 64.700 25.780 64.870 25.950 ;
        RECT 64.700 25.420 64.870 25.590 ;
        RECT 94.440 26.500 94.610 26.670 ;
        RECT 94.440 26.140 94.610 26.310 ;
        RECT 94.440 25.780 94.610 25.950 ;
        RECT 124.810 28.455 124.980 28.625 ;
        RECT 125.480 28.990 125.650 29.160 ;
        RECT 125.480 28.630 125.650 28.800 ;
        RECT 125.910 28.990 126.080 29.160 ;
        RECT 125.910 28.630 126.080 28.800 ;
        RECT 126.340 28.990 126.510 29.160 ;
        RECT 126.340 28.630 126.510 28.800 ;
        RECT 126.770 28.990 126.940 29.160 ;
        RECT 126.770 28.630 126.940 28.800 ;
        RECT 127.200 28.990 127.370 29.160 ;
        RECT 127.200 28.630 127.370 28.800 ;
        RECT 127.630 28.990 127.800 29.160 ;
        RECT 127.630 28.630 127.800 28.800 ;
        RECT 128.060 28.990 128.230 29.160 ;
        RECT 128.060 28.630 128.230 28.800 ;
        RECT 128.490 28.990 128.660 29.160 ;
        RECT 128.490 28.630 128.660 28.800 ;
        RECT 128.920 28.990 129.090 29.160 ;
        RECT 128.920 28.630 129.090 28.800 ;
        RECT 129.590 29.175 129.760 29.345 ;
        RECT 129.590 28.815 129.760 28.985 ;
        RECT 129.590 28.455 129.760 28.625 ;
        RECT 124.810 28.095 124.980 28.265 ;
        RECT 124.810 27.735 124.980 27.905 ;
        RECT 129.590 28.095 129.760 28.265 ;
        RECT 124.810 27.375 124.980 27.545 ;
        RECT 124.810 27.015 124.980 27.185 ;
        RECT 124.810 26.655 124.980 26.825 ;
        RECT 125.480 27.340 125.650 27.510 ;
        RECT 125.480 26.980 125.650 27.150 ;
        RECT 125.910 27.340 126.080 27.510 ;
        RECT 125.910 26.980 126.080 27.150 ;
        RECT 126.340 27.340 126.510 27.510 ;
        RECT 126.340 26.980 126.510 27.150 ;
        RECT 126.770 27.340 126.940 27.510 ;
        RECT 126.770 26.980 126.940 27.150 ;
        RECT 127.200 27.340 127.370 27.510 ;
        RECT 127.200 26.980 127.370 27.150 ;
        RECT 127.630 27.340 127.800 27.510 ;
        RECT 127.630 26.980 127.800 27.150 ;
        RECT 128.060 27.340 128.230 27.510 ;
        RECT 128.060 26.980 128.230 27.150 ;
        RECT 128.490 27.340 128.660 27.510 ;
        RECT 128.490 26.980 128.660 27.150 ;
        RECT 128.920 27.340 129.090 27.510 ;
        RECT 128.920 26.980 129.090 27.150 ;
        RECT 129.590 27.735 129.760 27.905 ;
        RECT 135.120 33.980 135.290 34.150 ;
        RECT 136.040 34.040 136.210 34.210 ;
        RECT 136.400 34.040 136.570 34.210 ;
        RECT 136.900 34.040 137.070 34.210 ;
        RECT 137.260 34.040 137.430 34.210 ;
        RECT 137.760 34.040 137.930 34.210 ;
        RECT 138.120 34.040 138.290 34.210 ;
        RECT 138.620 34.040 138.790 34.210 ;
        RECT 138.980 34.040 139.150 34.210 ;
        RECT 139.480 34.040 139.650 34.210 ;
        RECT 139.840 34.040 140.010 34.210 ;
        RECT 140.340 34.040 140.510 34.210 ;
        RECT 140.700 34.040 140.870 34.210 ;
        RECT 141.200 34.040 141.370 34.210 ;
        RECT 141.560 34.040 141.730 34.210 ;
        RECT 142.060 34.040 142.230 34.210 ;
        RECT 142.420 34.040 142.590 34.210 ;
        RECT 142.920 34.040 143.090 34.210 ;
        RECT 143.280 34.040 143.450 34.210 ;
        RECT 144.200 33.980 144.370 34.150 ;
        RECT 135.120 33.620 135.290 33.790 ;
        RECT 135.120 33.260 135.290 33.430 ;
        RECT 135.120 32.900 135.290 33.070 ;
        RECT 135.120 32.540 135.290 32.710 ;
        RECT 135.120 32.180 135.290 32.350 ;
        RECT 135.120 31.820 135.290 31.990 ;
        RECT 135.790 33.425 135.960 33.595 ;
        RECT 135.790 33.065 135.960 33.235 ;
        RECT 135.790 32.705 135.960 32.875 ;
        RECT 135.790 32.345 135.960 32.515 ;
        RECT 135.790 31.985 135.960 32.155 ;
        RECT 136.220 33.425 136.390 33.595 ;
        RECT 136.220 33.065 136.390 33.235 ;
        RECT 136.220 32.705 136.390 32.875 ;
        RECT 136.220 32.345 136.390 32.515 ;
        RECT 136.220 31.985 136.390 32.155 ;
        RECT 136.650 33.425 136.820 33.595 ;
        RECT 136.650 33.065 136.820 33.235 ;
        RECT 136.650 32.705 136.820 32.875 ;
        RECT 136.650 32.345 136.820 32.515 ;
        RECT 136.650 31.985 136.820 32.155 ;
        RECT 137.080 33.425 137.250 33.595 ;
        RECT 137.080 33.065 137.250 33.235 ;
        RECT 137.080 32.705 137.250 32.875 ;
        RECT 137.080 32.345 137.250 32.515 ;
        RECT 137.080 31.985 137.250 32.155 ;
        RECT 137.510 33.425 137.680 33.595 ;
        RECT 137.510 33.065 137.680 33.235 ;
        RECT 137.510 32.705 137.680 32.875 ;
        RECT 137.510 32.345 137.680 32.515 ;
        RECT 137.510 31.985 137.680 32.155 ;
        RECT 137.940 33.425 138.110 33.595 ;
        RECT 137.940 33.065 138.110 33.235 ;
        RECT 137.940 32.705 138.110 32.875 ;
        RECT 137.940 32.345 138.110 32.515 ;
        RECT 137.940 31.985 138.110 32.155 ;
        RECT 138.370 33.425 138.540 33.595 ;
        RECT 138.370 33.065 138.540 33.235 ;
        RECT 138.370 32.705 138.540 32.875 ;
        RECT 138.370 32.345 138.540 32.515 ;
        RECT 138.370 31.985 138.540 32.155 ;
        RECT 138.800 33.425 138.970 33.595 ;
        RECT 138.800 33.065 138.970 33.235 ;
        RECT 138.800 32.705 138.970 32.875 ;
        RECT 138.800 32.345 138.970 32.515 ;
        RECT 138.800 31.985 138.970 32.155 ;
        RECT 139.230 33.425 139.400 33.595 ;
        RECT 139.230 33.065 139.400 33.235 ;
        RECT 139.230 32.705 139.400 32.875 ;
        RECT 139.230 32.345 139.400 32.515 ;
        RECT 139.230 31.985 139.400 32.155 ;
        RECT 139.660 33.425 139.830 33.595 ;
        RECT 139.660 33.065 139.830 33.235 ;
        RECT 139.660 32.705 139.830 32.875 ;
        RECT 139.660 32.345 139.830 32.515 ;
        RECT 139.660 31.985 139.830 32.155 ;
        RECT 140.090 33.425 140.260 33.595 ;
        RECT 140.090 33.065 140.260 33.235 ;
        RECT 140.090 32.705 140.260 32.875 ;
        RECT 140.090 32.345 140.260 32.515 ;
        RECT 140.090 31.985 140.260 32.155 ;
        RECT 140.520 33.425 140.690 33.595 ;
        RECT 140.520 33.065 140.690 33.235 ;
        RECT 140.520 32.705 140.690 32.875 ;
        RECT 140.520 32.345 140.690 32.515 ;
        RECT 140.520 31.985 140.690 32.155 ;
        RECT 140.950 33.425 141.120 33.595 ;
        RECT 140.950 33.065 141.120 33.235 ;
        RECT 140.950 32.705 141.120 32.875 ;
        RECT 140.950 32.345 141.120 32.515 ;
        RECT 140.950 31.985 141.120 32.155 ;
        RECT 141.380 33.425 141.550 33.595 ;
        RECT 141.380 33.065 141.550 33.235 ;
        RECT 141.380 32.705 141.550 32.875 ;
        RECT 141.380 32.345 141.550 32.515 ;
        RECT 141.380 31.985 141.550 32.155 ;
        RECT 141.810 33.425 141.980 33.595 ;
        RECT 141.810 33.065 141.980 33.235 ;
        RECT 141.810 32.705 141.980 32.875 ;
        RECT 141.810 32.345 141.980 32.515 ;
        RECT 141.810 31.985 141.980 32.155 ;
        RECT 142.240 33.425 142.410 33.595 ;
        RECT 142.240 33.065 142.410 33.235 ;
        RECT 142.240 32.705 142.410 32.875 ;
        RECT 142.240 32.345 142.410 32.515 ;
        RECT 142.240 31.985 142.410 32.155 ;
        RECT 142.670 33.425 142.840 33.595 ;
        RECT 142.670 33.065 142.840 33.235 ;
        RECT 142.670 32.705 142.840 32.875 ;
        RECT 142.670 32.345 142.840 32.515 ;
        RECT 142.670 31.985 142.840 32.155 ;
        RECT 143.100 33.425 143.270 33.595 ;
        RECT 143.100 33.065 143.270 33.235 ;
        RECT 143.100 32.705 143.270 32.875 ;
        RECT 143.100 32.345 143.270 32.515 ;
        RECT 143.100 31.985 143.270 32.155 ;
        RECT 143.530 33.425 143.700 33.595 ;
        RECT 143.530 33.065 143.700 33.235 ;
        RECT 143.530 32.705 143.700 32.875 ;
        RECT 143.530 32.345 143.700 32.515 ;
        RECT 143.530 31.985 143.700 32.155 ;
        RECT 144.200 33.620 144.370 33.790 ;
        RECT 144.200 33.260 144.370 33.430 ;
        RECT 144.200 32.900 144.370 33.070 ;
        RECT 144.200 32.540 144.370 32.710 ;
        RECT 144.200 32.180 144.370 32.350 ;
        RECT 144.200 31.820 144.370 31.990 ;
        RECT 135.120 31.460 135.290 31.630 ;
        RECT 144.200 31.460 144.370 31.630 ;
        RECT 135.470 31.160 135.640 31.330 ;
        RECT 135.830 31.160 136.000 31.330 ;
        RECT 136.190 31.160 136.360 31.330 ;
        RECT 136.550 31.160 136.720 31.330 ;
        RECT 136.910 31.160 137.080 31.330 ;
        RECT 137.270 31.160 137.440 31.330 ;
        RECT 137.630 31.160 137.800 31.330 ;
        RECT 137.990 31.160 138.160 31.330 ;
        RECT 138.350 31.160 138.520 31.330 ;
        RECT 138.710 31.160 138.880 31.330 ;
        RECT 139.070 31.160 139.240 31.330 ;
        RECT 139.430 31.160 139.600 31.330 ;
        RECT 139.790 31.160 139.960 31.330 ;
        RECT 140.150 31.160 140.320 31.330 ;
        RECT 140.510 31.160 140.680 31.330 ;
        RECT 140.870 31.160 141.040 31.330 ;
        RECT 141.230 31.160 141.400 31.330 ;
        RECT 141.590 31.160 141.760 31.330 ;
        RECT 141.950 31.160 142.120 31.330 ;
        RECT 142.310 31.160 142.480 31.330 ;
        RECT 142.670 31.160 142.840 31.330 ;
        RECT 143.030 31.160 143.200 31.330 ;
        RECT 143.390 31.160 143.560 31.330 ;
        RECT 143.750 31.160 143.920 31.330 ;
        RECT 135.120 30.860 135.290 31.030 ;
        RECT 144.200 30.860 144.370 31.030 ;
        RECT 135.120 30.500 135.290 30.670 ;
        RECT 135.120 30.140 135.290 30.310 ;
        RECT 135.120 29.780 135.290 29.950 ;
        RECT 135.120 29.420 135.290 29.590 ;
        RECT 135.120 29.060 135.290 29.230 ;
        RECT 135.120 28.700 135.290 28.870 ;
        RECT 135.790 30.335 135.960 30.505 ;
        RECT 135.790 29.975 135.960 30.145 ;
        RECT 135.790 29.615 135.960 29.785 ;
        RECT 135.790 29.255 135.960 29.425 ;
        RECT 135.790 28.895 135.960 29.065 ;
        RECT 136.220 30.335 136.390 30.505 ;
        RECT 136.220 29.975 136.390 30.145 ;
        RECT 136.220 29.615 136.390 29.785 ;
        RECT 136.220 29.255 136.390 29.425 ;
        RECT 136.220 28.895 136.390 29.065 ;
        RECT 136.650 30.335 136.820 30.505 ;
        RECT 136.650 29.975 136.820 30.145 ;
        RECT 136.650 29.615 136.820 29.785 ;
        RECT 136.650 29.255 136.820 29.425 ;
        RECT 136.650 28.895 136.820 29.065 ;
        RECT 137.080 30.335 137.250 30.505 ;
        RECT 137.080 29.975 137.250 30.145 ;
        RECT 137.080 29.615 137.250 29.785 ;
        RECT 137.080 29.255 137.250 29.425 ;
        RECT 137.080 28.895 137.250 29.065 ;
        RECT 137.510 30.335 137.680 30.505 ;
        RECT 137.510 29.975 137.680 30.145 ;
        RECT 137.510 29.615 137.680 29.785 ;
        RECT 137.510 29.255 137.680 29.425 ;
        RECT 137.510 28.895 137.680 29.065 ;
        RECT 137.940 30.335 138.110 30.505 ;
        RECT 137.940 29.975 138.110 30.145 ;
        RECT 137.940 29.615 138.110 29.785 ;
        RECT 137.940 29.255 138.110 29.425 ;
        RECT 137.940 28.895 138.110 29.065 ;
        RECT 138.370 30.335 138.540 30.505 ;
        RECT 138.370 29.975 138.540 30.145 ;
        RECT 138.370 29.615 138.540 29.785 ;
        RECT 138.370 29.255 138.540 29.425 ;
        RECT 138.370 28.895 138.540 29.065 ;
        RECT 138.800 30.335 138.970 30.505 ;
        RECT 138.800 29.975 138.970 30.145 ;
        RECT 138.800 29.615 138.970 29.785 ;
        RECT 138.800 29.255 138.970 29.425 ;
        RECT 138.800 28.895 138.970 29.065 ;
        RECT 139.230 30.335 139.400 30.505 ;
        RECT 139.230 29.975 139.400 30.145 ;
        RECT 139.230 29.615 139.400 29.785 ;
        RECT 139.230 29.255 139.400 29.425 ;
        RECT 139.230 28.895 139.400 29.065 ;
        RECT 139.660 30.335 139.830 30.505 ;
        RECT 139.660 29.975 139.830 30.145 ;
        RECT 139.660 29.615 139.830 29.785 ;
        RECT 139.660 29.255 139.830 29.425 ;
        RECT 139.660 28.895 139.830 29.065 ;
        RECT 140.090 30.335 140.260 30.505 ;
        RECT 140.090 29.975 140.260 30.145 ;
        RECT 140.090 29.615 140.260 29.785 ;
        RECT 140.090 29.255 140.260 29.425 ;
        RECT 140.090 28.895 140.260 29.065 ;
        RECT 140.520 30.335 140.690 30.505 ;
        RECT 140.520 29.975 140.690 30.145 ;
        RECT 140.520 29.615 140.690 29.785 ;
        RECT 140.520 29.255 140.690 29.425 ;
        RECT 140.520 28.895 140.690 29.065 ;
        RECT 140.950 30.335 141.120 30.505 ;
        RECT 140.950 29.975 141.120 30.145 ;
        RECT 140.950 29.615 141.120 29.785 ;
        RECT 140.950 29.255 141.120 29.425 ;
        RECT 140.950 28.895 141.120 29.065 ;
        RECT 141.380 30.335 141.550 30.505 ;
        RECT 141.380 29.975 141.550 30.145 ;
        RECT 141.380 29.615 141.550 29.785 ;
        RECT 141.380 29.255 141.550 29.425 ;
        RECT 141.380 28.895 141.550 29.065 ;
        RECT 141.810 30.335 141.980 30.505 ;
        RECT 141.810 29.975 141.980 30.145 ;
        RECT 141.810 29.615 141.980 29.785 ;
        RECT 141.810 29.255 141.980 29.425 ;
        RECT 141.810 28.895 141.980 29.065 ;
        RECT 142.240 30.335 142.410 30.505 ;
        RECT 142.240 29.975 142.410 30.145 ;
        RECT 142.240 29.615 142.410 29.785 ;
        RECT 142.240 29.255 142.410 29.425 ;
        RECT 142.240 28.895 142.410 29.065 ;
        RECT 142.670 30.335 142.840 30.505 ;
        RECT 142.670 29.975 142.840 30.145 ;
        RECT 142.670 29.615 142.840 29.785 ;
        RECT 142.670 29.255 142.840 29.425 ;
        RECT 142.670 28.895 142.840 29.065 ;
        RECT 143.100 30.335 143.270 30.505 ;
        RECT 143.100 29.975 143.270 30.145 ;
        RECT 143.100 29.615 143.270 29.785 ;
        RECT 143.100 29.255 143.270 29.425 ;
        RECT 143.100 28.895 143.270 29.065 ;
        RECT 143.530 30.335 143.700 30.505 ;
        RECT 143.530 29.975 143.700 30.145 ;
        RECT 143.530 29.615 143.700 29.785 ;
        RECT 143.530 29.255 143.700 29.425 ;
        RECT 143.530 28.895 143.700 29.065 ;
        RECT 144.200 30.500 144.370 30.670 ;
        RECT 144.200 30.140 144.370 30.310 ;
        RECT 144.200 29.780 144.370 29.950 ;
        RECT 144.200 29.420 144.370 29.590 ;
        RECT 144.200 29.060 144.370 29.230 ;
        RECT 144.200 28.700 144.370 28.870 ;
        RECT 135.120 28.340 135.290 28.510 ;
        RECT 136.040 28.280 136.210 28.450 ;
        RECT 136.400 28.280 136.570 28.450 ;
        RECT 136.900 28.280 137.070 28.450 ;
        RECT 137.260 28.280 137.430 28.450 ;
        RECT 137.760 28.280 137.930 28.450 ;
        RECT 138.120 28.280 138.290 28.450 ;
        RECT 138.620 28.280 138.790 28.450 ;
        RECT 138.980 28.280 139.150 28.450 ;
        RECT 139.480 28.280 139.650 28.450 ;
        RECT 139.840 28.280 140.010 28.450 ;
        RECT 140.340 28.280 140.510 28.450 ;
        RECT 140.700 28.280 140.870 28.450 ;
        RECT 141.200 28.280 141.370 28.450 ;
        RECT 141.560 28.280 141.730 28.450 ;
        RECT 142.060 28.280 142.230 28.450 ;
        RECT 142.420 28.280 142.590 28.450 ;
        RECT 142.920 28.280 143.090 28.450 ;
        RECT 143.280 28.280 143.450 28.450 ;
        RECT 144.200 28.340 144.370 28.510 ;
        RECT 129.590 27.375 129.760 27.545 ;
        RECT 129.590 27.015 129.760 27.185 ;
        RECT 129.590 26.655 129.760 26.825 ;
        RECT 124.810 26.295 124.980 26.465 ;
        RECT 125.730 26.325 125.900 26.495 ;
        RECT 126.090 26.325 126.260 26.495 ;
        RECT 126.590 26.325 126.760 26.495 ;
        RECT 126.950 26.325 127.120 26.495 ;
        RECT 127.450 26.325 127.620 26.495 ;
        RECT 127.810 26.325 127.980 26.495 ;
        RECT 128.310 26.325 128.480 26.495 ;
        RECT 128.670 26.325 128.840 26.495 ;
        RECT 129.590 26.295 129.760 26.465 ;
        RECT 135.120 26.845 135.290 27.015 ;
        RECT 135.120 26.485 135.290 26.655 ;
        RECT 136.040 26.600 136.210 26.770 ;
        RECT 136.400 26.600 136.570 26.770 ;
        RECT 136.900 26.600 137.070 26.770 ;
        RECT 137.260 26.600 137.430 26.770 ;
        RECT 137.760 26.600 137.930 26.770 ;
        RECT 138.120 26.600 138.290 26.770 ;
        RECT 138.620 26.600 138.790 26.770 ;
        RECT 138.980 26.600 139.150 26.770 ;
        RECT 139.480 26.600 139.650 26.770 ;
        RECT 139.840 26.600 140.010 26.770 ;
        RECT 140.340 26.600 140.510 26.770 ;
        RECT 140.700 26.600 140.870 26.770 ;
        RECT 141.200 26.600 141.370 26.770 ;
        RECT 141.560 26.600 141.730 26.770 ;
        RECT 142.060 26.600 142.230 26.770 ;
        RECT 142.420 26.600 142.590 26.770 ;
        RECT 142.920 26.600 143.090 26.770 ;
        RECT 143.280 26.600 143.450 26.770 ;
        RECT 144.200 26.845 144.370 27.015 ;
        RECT 144.200 26.485 144.370 26.655 ;
        RECT 135.120 26.125 135.290 26.295 ;
        RECT 65.715 25.310 65.885 25.480 ;
        RECT 66.075 25.310 66.245 25.480 ;
        RECT 66.435 25.310 66.605 25.480 ;
        RECT 66.795 25.310 66.965 25.480 ;
        RECT 67.155 25.310 67.325 25.480 ;
        RECT 67.515 25.310 67.685 25.480 ;
        RECT 68.310 25.310 68.480 25.480 ;
        RECT 68.670 25.310 68.840 25.480 ;
        RECT 69.030 25.310 69.200 25.480 ;
        RECT 69.390 25.310 69.560 25.480 ;
        RECT 69.750 25.310 69.920 25.480 ;
        RECT 70.590 25.310 70.760 25.480 ;
        RECT 70.950 25.310 71.120 25.480 ;
        RECT 71.310 25.310 71.480 25.480 ;
        RECT 71.670 25.310 71.840 25.480 ;
        RECT 72.030 25.310 72.200 25.480 ;
        RECT 72.870 25.310 73.040 25.480 ;
        RECT 73.230 25.310 73.400 25.480 ;
        RECT 73.590 25.310 73.760 25.480 ;
        RECT 73.950 25.310 74.120 25.480 ;
        RECT 74.310 25.310 74.480 25.480 ;
        RECT 75.150 25.310 75.320 25.480 ;
        RECT 75.510 25.310 75.680 25.480 ;
        RECT 75.870 25.310 76.040 25.480 ;
        RECT 76.230 25.310 76.400 25.480 ;
        RECT 76.590 25.310 76.760 25.480 ;
        RECT 77.395 25.310 77.565 25.480 ;
        RECT 77.755 25.310 77.925 25.480 ;
        RECT 78.115 25.310 78.285 25.480 ;
        RECT 78.475 25.310 78.645 25.480 ;
        RECT 78.835 25.310 79.005 25.480 ;
        RECT 79.195 25.310 79.365 25.480 ;
        RECT 79.955 25.310 80.125 25.480 ;
        RECT 80.315 25.310 80.485 25.480 ;
        RECT 80.675 25.310 80.845 25.480 ;
        RECT 81.035 25.310 81.205 25.480 ;
        RECT 81.395 25.310 81.565 25.480 ;
        RECT 81.755 25.310 81.925 25.480 ;
        RECT 82.550 25.310 82.720 25.480 ;
        RECT 82.910 25.310 83.080 25.480 ;
        RECT 83.270 25.310 83.440 25.480 ;
        RECT 83.630 25.310 83.800 25.480 ;
        RECT 83.990 25.310 84.160 25.480 ;
        RECT 84.830 25.310 85.000 25.480 ;
        RECT 85.190 25.310 85.360 25.480 ;
        RECT 85.550 25.310 85.720 25.480 ;
        RECT 85.910 25.310 86.080 25.480 ;
        RECT 86.270 25.310 86.440 25.480 ;
        RECT 87.110 25.310 87.280 25.480 ;
        RECT 87.470 25.310 87.640 25.480 ;
        RECT 87.830 25.310 88.000 25.480 ;
        RECT 88.190 25.310 88.360 25.480 ;
        RECT 88.550 25.310 88.720 25.480 ;
        RECT 89.390 25.310 89.560 25.480 ;
        RECT 89.750 25.310 89.920 25.480 ;
        RECT 90.110 25.310 90.280 25.480 ;
        RECT 90.470 25.310 90.640 25.480 ;
        RECT 90.830 25.310 91.000 25.480 ;
        RECT 91.635 25.310 91.805 25.480 ;
        RECT 91.995 25.310 92.165 25.480 ;
        RECT 92.355 25.310 92.525 25.480 ;
        RECT 92.715 25.310 92.885 25.480 ;
        RECT 93.075 25.310 93.245 25.480 ;
        RECT 93.435 25.310 93.605 25.480 ;
        RECT 94.440 25.420 94.610 25.590 ;
        RECT 135.120 25.765 135.290 25.935 ;
        RECT 135.120 25.405 135.290 25.575 ;
        RECT 64.700 25.060 64.870 25.230 ;
        RECT 94.440 25.060 94.610 25.230 ;
        RECT 64.700 24.700 64.870 24.870 ;
        RECT 65.330 24.725 65.500 24.895 ;
        RECT 66.610 24.725 66.780 24.895 ;
        RECT 67.890 24.725 68.060 24.895 ;
        RECT 70.170 24.725 70.340 24.895 ;
        RECT 72.450 24.725 72.620 24.895 ;
        RECT 74.730 24.725 74.900 24.895 ;
        RECT 77.010 24.725 77.180 24.895 ;
        RECT 78.290 24.725 78.460 24.895 ;
        RECT 79.570 24.725 79.740 24.895 ;
        RECT 80.850 24.725 81.020 24.895 ;
        RECT 82.130 24.725 82.300 24.895 ;
        RECT 84.410 24.725 84.580 24.895 ;
        RECT 86.690 24.725 86.860 24.895 ;
        RECT 88.970 24.725 89.140 24.895 ;
        RECT 91.250 24.725 91.420 24.895 ;
        RECT 92.530 24.725 92.700 24.895 ;
        RECT 93.810 24.725 93.980 24.895 ;
        RECT 94.440 24.700 94.610 24.870 ;
        RECT 64.700 24.340 64.870 24.510 ;
        RECT 64.700 23.980 64.870 24.150 ;
        RECT 68.310 24.140 68.480 24.310 ;
        RECT 68.670 24.140 68.840 24.310 ;
        RECT 69.030 24.140 69.200 24.310 ;
        RECT 69.390 24.140 69.560 24.310 ;
        RECT 69.750 24.140 69.920 24.310 ;
        RECT 70.590 24.140 70.760 24.310 ;
        RECT 70.950 24.140 71.120 24.310 ;
        RECT 71.310 24.140 71.480 24.310 ;
        RECT 71.670 24.140 71.840 24.310 ;
        RECT 72.030 24.140 72.200 24.310 ;
        RECT 72.870 24.140 73.040 24.310 ;
        RECT 73.230 24.140 73.400 24.310 ;
        RECT 73.590 24.140 73.760 24.310 ;
        RECT 73.950 24.140 74.120 24.310 ;
        RECT 74.310 24.140 74.480 24.310 ;
        RECT 75.150 24.140 75.320 24.310 ;
        RECT 75.510 24.140 75.680 24.310 ;
        RECT 75.870 24.140 76.040 24.310 ;
        RECT 76.230 24.140 76.400 24.310 ;
        RECT 76.590 24.140 76.760 24.310 ;
        RECT 77.395 24.140 77.565 24.310 ;
        RECT 77.755 24.140 77.925 24.310 ;
        RECT 78.115 24.140 78.285 24.310 ;
        RECT 78.475 24.140 78.645 24.310 ;
        RECT 78.835 24.140 79.005 24.310 ;
        RECT 79.195 24.140 79.365 24.310 ;
        RECT 79.955 24.140 80.125 24.310 ;
        RECT 80.315 24.140 80.485 24.310 ;
        RECT 80.675 24.140 80.845 24.310 ;
        RECT 81.035 24.140 81.205 24.310 ;
        RECT 81.395 24.140 81.565 24.310 ;
        RECT 81.755 24.140 81.925 24.310 ;
        RECT 82.550 24.140 82.720 24.310 ;
        RECT 82.910 24.140 83.080 24.310 ;
        RECT 83.270 24.140 83.440 24.310 ;
        RECT 83.630 24.140 83.800 24.310 ;
        RECT 83.990 24.140 84.160 24.310 ;
        RECT 84.830 24.140 85.000 24.310 ;
        RECT 85.190 24.140 85.360 24.310 ;
        RECT 85.550 24.140 85.720 24.310 ;
        RECT 85.910 24.140 86.080 24.310 ;
        RECT 86.270 24.140 86.440 24.310 ;
        RECT 87.110 24.140 87.280 24.310 ;
        RECT 87.470 24.140 87.640 24.310 ;
        RECT 87.830 24.140 88.000 24.310 ;
        RECT 88.190 24.140 88.360 24.310 ;
        RECT 88.550 24.140 88.720 24.310 ;
        RECT 89.390 24.140 89.560 24.310 ;
        RECT 89.750 24.140 89.920 24.310 ;
        RECT 90.110 24.140 90.280 24.310 ;
        RECT 90.470 24.140 90.640 24.310 ;
        RECT 90.830 24.140 91.000 24.310 ;
        RECT 94.440 24.340 94.610 24.510 ;
        RECT 94.440 23.980 94.610 24.150 ;
        RECT 65.050 23.590 65.220 23.760 ;
        RECT 65.410 23.590 65.580 23.760 ;
        RECT 65.770 23.590 65.940 23.760 ;
        RECT 66.130 23.590 66.300 23.760 ;
        RECT 66.490 23.590 66.660 23.760 ;
        RECT 66.850 23.590 67.020 23.760 ;
        RECT 67.210 23.590 67.380 23.760 ;
        RECT 67.570 23.590 67.740 23.760 ;
        RECT 67.930 23.590 68.100 23.760 ;
        RECT 68.290 23.590 68.460 23.760 ;
        RECT 68.650 23.590 68.820 23.760 ;
        RECT 69.010 23.590 69.180 23.760 ;
        RECT 69.370 23.590 69.540 23.760 ;
        RECT 69.730 23.590 69.900 23.760 ;
        RECT 70.090 23.590 70.260 23.760 ;
        RECT 70.450 23.590 70.620 23.760 ;
        RECT 70.810 23.590 70.980 23.760 ;
        RECT 71.170 23.590 71.340 23.760 ;
        RECT 71.530 23.590 71.700 23.760 ;
        RECT 71.890 23.590 72.060 23.760 ;
        RECT 72.250 23.590 72.420 23.760 ;
        RECT 72.610 23.590 72.780 23.760 ;
        RECT 72.970 23.590 73.140 23.760 ;
        RECT 73.330 23.590 73.500 23.760 ;
        RECT 73.690 23.590 73.860 23.760 ;
        RECT 74.050 23.590 74.220 23.760 ;
        RECT 74.410 23.590 74.580 23.760 ;
        RECT 74.770 23.590 74.940 23.760 ;
        RECT 75.130 23.590 75.300 23.760 ;
        RECT 75.490 23.590 75.660 23.760 ;
        RECT 75.850 23.590 76.020 23.760 ;
        RECT 76.210 23.590 76.380 23.760 ;
        RECT 76.570 23.590 76.740 23.760 ;
        RECT 76.930 23.590 77.100 23.760 ;
        RECT 77.290 23.590 77.460 23.760 ;
        RECT 77.650 23.590 77.820 23.760 ;
        RECT 78.010 23.590 78.180 23.760 ;
        RECT 78.370 23.590 78.540 23.760 ;
        RECT 78.730 23.590 78.900 23.760 ;
        RECT 79.090 23.590 79.260 23.760 ;
        RECT 79.450 23.590 79.620 23.760 ;
        RECT 79.810 23.590 79.980 23.760 ;
        RECT 80.170 23.590 80.340 23.760 ;
        RECT 80.530 23.590 80.700 23.760 ;
        RECT 80.890 23.590 81.060 23.760 ;
        RECT 81.250 23.590 81.420 23.760 ;
        RECT 81.610 23.590 81.780 23.760 ;
        RECT 81.970 23.590 82.140 23.760 ;
        RECT 82.330 23.590 82.500 23.760 ;
        RECT 82.690 23.590 82.860 23.760 ;
        RECT 83.050 23.590 83.220 23.760 ;
        RECT 83.410 23.590 83.580 23.760 ;
        RECT 83.770 23.590 83.940 23.760 ;
        RECT 84.130 23.590 84.300 23.760 ;
        RECT 84.490 23.590 84.660 23.760 ;
        RECT 84.850 23.590 85.020 23.760 ;
        RECT 85.210 23.590 85.380 23.760 ;
        RECT 85.570 23.590 85.740 23.760 ;
        RECT 85.930 23.590 86.100 23.760 ;
        RECT 86.290 23.590 86.460 23.760 ;
        RECT 86.650 23.590 86.820 23.760 ;
        RECT 87.010 23.590 87.180 23.760 ;
        RECT 87.370 23.590 87.540 23.760 ;
        RECT 87.730 23.590 87.900 23.760 ;
        RECT 88.090 23.590 88.260 23.760 ;
        RECT 88.450 23.590 88.620 23.760 ;
        RECT 88.810 23.590 88.980 23.760 ;
        RECT 89.170 23.590 89.340 23.760 ;
        RECT 89.530 23.590 89.700 23.760 ;
        RECT 89.890 23.590 90.060 23.760 ;
        RECT 90.250 23.590 90.420 23.760 ;
        RECT 90.610 23.590 90.780 23.760 ;
        RECT 90.970 23.590 91.140 23.760 ;
        RECT 91.330 23.590 91.500 23.760 ;
        RECT 91.690 23.590 91.860 23.760 ;
        RECT 92.050 23.590 92.220 23.760 ;
        RECT 92.410 23.590 92.580 23.760 ;
        RECT 92.770 23.590 92.940 23.760 ;
        RECT 93.130 23.590 93.300 23.760 ;
        RECT 93.490 23.590 93.660 23.760 ;
        RECT 93.850 23.590 94.020 23.760 ;
        RECT 124.810 24.575 124.980 24.745 ;
        RECT 125.730 24.695 125.900 24.865 ;
        RECT 126.090 24.695 126.260 24.865 ;
        RECT 126.590 24.695 126.760 24.865 ;
        RECT 126.950 24.695 127.120 24.865 ;
        RECT 127.450 24.695 127.620 24.865 ;
        RECT 127.810 24.695 127.980 24.865 ;
        RECT 128.310 24.695 128.480 24.865 ;
        RECT 128.670 24.695 128.840 24.865 ;
        RECT 135.790 25.945 135.960 26.115 ;
        RECT 135.790 25.585 135.960 25.755 ;
        RECT 136.220 25.945 136.390 26.115 ;
        RECT 136.220 25.585 136.390 25.755 ;
        RECT 136.650 25.945 136.820 26.115 ;
        RECT 136.650 25.585 136.820 25.755 ;
        RECT 137.080 25.945 137.250 26.115 ;
        RECT 137.080 25.585 137.250 25.755 ;
        RECT 137.510 25.945 137.680 26.115 ;
        RECT 137.510 25.585 137.680 25.755 ;
        RECT 137.940 25.945 138.110 26.115 ;
        RECT 137.940 25.585 138.110 25.755 ;
        RECT 138.370 25.945 138.540 26.115 ;
        RECT 138.370 25.585 138.540 25.755 ;
        RECT 138.800 25.945 138.970 26.115 ;
        RECT 138.800 25.585 138.970 25.755 ;
        RECT 139.230 25.945 139.400 26.115 ;
        RECT 139.230 25.585 139.400 25.755 ;
        RECT 139.660 25.945 139.830 26.115 ;
        RECT 139.660 25.585 139.830 25.755 ;
        RECT 140.090 25.945 140.260 26.115 ;
        RECT 140.090 25.585 140.260 25.755 ;
        RECT 140.520 25.945 140.690 26.115 ;
        RECT 140.520 25.585 140.690 25.755 ;
        RECT 140.950 25.945 141.120 26.115 ;
        RECT 140.950 25.585 141.120 25.755 ;
        RECT 141.380 25.945 141.550 26.115 ;
        RECT 141.380 25.585 141.550 25.755 ;
        RECT 141.810 25.945 141.980 26.115 ;
        RECT 141.810 25.585 141.980 25.755 ;
        RECT 142.240 25.945 142.410 26.115 ;
        RECT 142.240 25.585 142.410 25.755 ;
        RECT 142.670 25.945 142.840 26.115 ;
        RECT 142.670 25.585 142.840 25.755 ;
        RECT 143.100 25.945 143.270 26.115 ;
        RECT 143.100 25.585 143.270 25.755 ;
        RECT 143.530 25.945 143.700 26.115 ;
        RECT 143.530 25.585 143.700 25.755 ;
        RECT 144.200 26.125 144.370 26.295 ;
        RECT 144.200 25.765 144.370 25.935 ;
        RECT 144.200 25.405 144.370 25.575 ;
        RECT 135.120 25.045 135.290 25.215 ;
        RECT 144.200 25.045 144.370 25.215 ;
        RECT 135.470 24.745 135.640 24.915 ;
        RECT 135.830 24.745 136.000 24.915 ;
        RECT 136.190 24.745 136.360 24.915 ;
        RECT 136.550 24.745 136.720 24.915 ;
        RECT 136.910 24.745 137.080 24.915 ;
        RECT 137.270 24.745 137.440 24.915 ;
        RECT 137.630 24.745 137.800 24.915 ;
        RECT 137.990 24.745 138.160 24.915 ;
        RECT 138.350 24.745 138.520 24.915 ;
        RECT 138.710 24.745 138.880 24.915 ;
        RECT 139.070 24.745 139.240 24.915 ;
        RECT 139.430 24.745 139.600 24.915 ;
        RECT 139.790 24.745 139.960 24.915 ;
        RECT 140.150 24.745 140.320 24.915 ;
        RECT 140.510 24.745 140.680 24.915 ;
        RECT 140.870 24.745 141.040 24.915 ;
        RECT 141.230 24.745 141.400 24.915 ;
        RECT 141.590 24.745 141.760 24.915 ;
        RECT 141.950 24.745 142.120 24.915 ;
        RECT 142.310 24.745 142.480 24.915 ;
        RECT 142.670 24.745 142.840 24.915 ;
        RECT 143.030 24.745 143.200 24.915 ;
        RECT 143.390 24.745 143.560 24.915 ;
        RECT 143.750 24.745 143.920 24.915 ;
        RECT 129.590 24.575 129.760 24.745 ;
        RECT 124.810 24.215 124.980 24.385 ;
        RECT 124.810 23.855 124.980 24.025 ;
        RECT 124.810 23.495 124.980 23.665 ;
        RECT 125.480 24.040 125.650 24.210 ;
        RECT 125.480 23.680 125.650 23.850 ;
        RECT 125.910 24.040 126.080 24.210 ;
        RECT 125.910 23.680 126.080 23.850 ;
        RECT 126.340 24.040 126.510 24.210 ;
        RECT 126.340 23.680 126.510 23.850 ;
        RECT 126.770 24.040 126.940 24.210 ;
        RECT 126.770 23.680 126.940 23.850 ;
        RECT 127.200 24.040 127.370 24.210 ;
        RECT 127.200 23.680 127.370 23.850 ;
        RECT 127.630 24.040 127.800 24.210 ;
        RECT 127.630 23.680 127.800 23.850 ;
        RECT 128.060 24.040 128.230 24.210 ;
        RECT 128.060 23.680 128.230 23.850 ;
        RECT 128.490 24.040 128.660 24.210 ;
        RECT 128.490 23.680 128.660 23.850 ;
        RECT 128.920 24.040 129.090 24.210 ;
        RECT 128.920 23.680 129.090 23.850 ;
        RECT 129.590 24.215 129.760 24.385 ;
        RECT 129.590 23.855 129.760 24.025 ;
        RECT 129.590 23.495 129.760 23.665 ;
        RECT 124.810 23.135 124.980 23.305 ;
        RECT 125.730 23.025 125.900 23.195 ;
        RECT 126.090 23.025 126.260 23.195 ;
        RECT 126.590 23.025 126.760 23.195 ;
        RECT 126.950 23.025 127.120 23.195 ;
        RECT 127.450 23.025 127.620 23.195 ;
        RECT 127.810 23.025 127.980 23.195 ;
        RECT 128.310 23.025 128.480 23.195 ;
        RECT 128.670 23.025 128.840 23.195 ;
        RECT 129.590 23.135 129.760 23.305 ;
        RECT 124.810 22.775 124.980 22.945 ;
        RECT 129.590 22.775 129.760 22.945 ;
        RECT 125.160 22.475 125.330 22.645 ;
        RECT 125.520 22.475 125.690 22.645 ;
        RECT 125.880 22.475 126.050 22.645 ;
        RECT 126.240 22.475 126.410 22.645 ;
        RECT 126.600 22.475 126.770 22.645 ;
        RECT 126.960 22.475 127.130 22.645 ;
        RECT 127.320 22.475 127.490 22.645 ;
        RECT 127.680 22.475 127.850 22.645 ;
        RECT 128.040 22.475 128.210 22.645 ;
        RECT 128.400 22.475 128.570 22.645 ;
        RECT 128.760 22.475 128.930 22.645 ;
        RECT 129.120 22.475 129.290 22.645 ;
        RECT 135.470 22.140 135.640 22.310 ;
        RECT 135.830 22.140 136.000 22.310 ;
        RECT 136.190 22.140 136.360 22.310 ;
        RECT 136.550 22.140 136.720 22.310 ;
        RECT 136.910 22.140 137.080 22.310 ;
        RECT 137.270 22.140 137.440 22.310 ;
        RECT 137.630 22.140 137.800 22.310 ;
        RECT 137.990 22.140 138.160 22.310 ;
        RECT 138.350 22.140 138.520 22.310 ;
        RECT 138.710 22.140 138.880 22.310 ;
        RECT 139.070 22.140 139.240 22.310 ;
        RECT 139.430 22.140 139.600 22.310 ;
        RECT 139.790 22.140 139.960 22.310 ;
        RECT 140.150 22.140 140.320 22.310 ;
        RECT 140.510 22.140 140.680 22.310 ;
        RECT 140.870 22.140 141.040 22.310 ;
        RECT 141.230 22.140 141.400 22.310 ;
        RECT 141.590 22.140 141.760 22.310 ;
        RECT 141.950 22.140 142.120 22.310 ;
        RECT 142.310 22.140 142.480 22.310 ;
        RECT 142.670 22.140 142.840 22.310 ;
        RECT 143.030 22.140 143.200 22.310 ;
        RECT 143.390 22.140 143.560 22.310 ;
        RECT 143.750 22.140 143.920 22.310 ;
        RECT 69.540 21.960 69.710 22.130 ;
        RECT 69.900 21.960 70.070 22.130 ;
        RECT 70.260 21.960 70.430 22.130 ;
        RECT 70.620 21.960 70.790 22.130 ;
        RECT 70.980 21.960 71.150 22.130 ;
        RECT 71.340 21.960 71.510 22.130 ;
        RECT 71.700 21.960 71.870 22.130 ;
        RECT 72.060 21.960 72.230 22.130 ;
        RECT 72.420 21.960 72.590 22.130 ;
        RECT 72.780 21.960 72.950 22.130 ;
        RECT 73.140 21.960 73.310 22.130 ;
        RECT 73.500 21.960 73.670 22.130 ;
        RECT 73.860 21.960 74.030 22.130 ;
        RECT 74.220 21.960 74.390 22.130 ;
        RECT 74.580 21.960 74.750 22.130 ;
        RECT 74.940 21.960 75.110 22.130 ;
        RECT 75.300 21.960 75.470 22.130 ;
        RECT 75.660 21.960 75.830 22.130 ;
        RECT 76.020 21.960 76.190 22.130 ;
        RECT 76.380 21.960 76.550 22.130 ;
        RECT 76.740 21.960 76.910 22.130 ;
        RECT 77.100 21.960 77.270 22.130 ;
        RECT 77.460 21.960 77.630 22.130 ;
        RECT 77.820 21.960 77.990 22.130 ;
        RECT 78.180 21.960 78.350 22.130 ;
        RECT 78.540 21.960 78.710 22.130 ;
        RECT 78.900 21.960 79.070 22.130 ;
        RECT 79.260 21.960 79.430 22.130 ;
        RECT 79.620 21.960 79.790 22.130 ;
        RECT 79.980 21.960 80.150 22.130 ;
        RECT 80.340 21.960 80.510 22.130 ;
        RECT 80.700 21.960 80.870 22.130 ;
        RECT 81.060 21.960 81.230 22.130 ;
        RECT 81.420 21.960 81.590 22.130 ;
        RECT 81.780 21.960 81.950 22.130 ;
        RECT 82.140 21.960 82.310 22.130 ;
        RECT 82.500 21.960 82.670 22.130 ;
        RECT 82.860 21.960 83.030 22.130 ;
        RECT 83.220 21.960 83.390 22.130 ;
        RECT 83.580 21.960 83.750 22.130 ;
        RECT 83.940 21.960 84.110 22.130 ;
        RECT 84.300 21.960 84.470 22.130 ;
        RECT 84.660 21.960 84.830 22.130 ;
        RECT 85.020 21.960 85.190 22.130 ;
        RECT 85.380 21.960 85.550 22.130 ;
        RECT 85.740 21.960 85.910 22.130 ;
        RECT 86.100 21.960 86.270 22.130 ;
        RECT 86.460 21.960 86.630 22.130 ;
        RECT 86.820 21.960 86.990 22.130 ;
        RECT 87.180 21.960 87.350 22.130 ;
        RECT 87.540 21.960 87.710 22.130 ;
        RECT 87.900 21.960 88.070 22.130 ;
        RECT 88.260 21.960 88.430 22.130 ;
        RECT 88.620 21.960 88.790 22.130 ;
        RECT 88.980 21.960 89.150 22.130 ;
        RECT 89.340 21.960 89.510 22.130 ;
        RECT 69.190 21.660 69.360 21.830 ;
        RECT 89.890 21.660 90.060 21.830 ;
        RECT 69.190 21.300 69.360 21.470 ;
        RECT 70.245 21.410 70.415 21.580 ;
        RECT 70.605 21.410 70.775 21.580 ;
        RECT 70.965 21.410 71.135 21.580 ;
        RECT 71.325 21.410 71.495 21.580 ;
        RECT 71.685 21.410 71.855 21.580 ;
        RECT 72.045 21.410 72.215 21.580 ;
        RECT 72.840 21.410 73.010 21.580 ;
        RECT 73.200 21.410 73.370 21.580 ;
        RECT 73.560 21.410 73.730 21.580 ;
        RECT 73.920 21.410 74.090 21.580 ;
        RECT 74.280 21.410 74.450 21.580 ;
        RECT 75.120 21.410 75.290 21.580 ;
        RECT 75.480 21.410 75.650 21.580 ;
        RECT 75.840 21.410 76.010 21.580 ;
        RECT 76.200 21.410 76.370 21.580 ;
        RECT 76.560 21.410 76.730 21.580 ;
        RECT 77.365 21.410 77.535 21.580 ;
        RECT 77.725 21.410 77.895 21.580 ;
        RECT 78.085 21.410 78.255 21.580 ;
        RECT 78.445 21.410 78.615 21.580 ;
        RECT 78.805 21.410 78.975 21.580 ;
        RECT 79.165 21.410 79.335 21.580 ;
        RECT 79.925 21.410 80.095 21.580 ;
        RECT 80.285 21.410 80.455 21.580 ;
        RECT 80.645 21.410 80.815 21.580 ;
        RECT 81.005 21.410 81.175 21.580 ;
        RECT 81.365 21.410 81.535 21.580 ;
        RECT 81.725 21.410 81.895 21.580 ;
        RECT 82.520 21.410 82.690 21.580 ;
        RECT 82.880 21.410 83.050 21.580 ;
        RECT 83.240 21.410 83.410 21.580 ;
        RECT 83.600 21.410 83.770 21.580 ;
        RECT 83.960 21.410 84.130 21.580 ;
        RECT 84.800 21.410 84.970 21.580 ;
        RECT 85.160 21.410 85.330 21.580 ;
        RECT 85.520 21.410 85.690 21.580 ;
        RECT 85.880 21.410 86.050 21.580 ;
        RECT 86.240 21.410 86.410 21.580 ;
        RECT 87.045 21.410 87.215 21.580 ;
        RECT 87.405 21.410 87.575 21.580 ;
        RECT 87.765 21.410 87.935 21.580 ;
        RECT 88.125 21.410 88.295 21.580 ;
        RECT 88.485 21.410 88.655 21.580 ;
        RECT 88.845 21.410 89.015 21.580 ;
        RECT 89.890 21.300 90.060 21.470 ;
        RECT 69.190 20.940 69.360 21.110 ;
        RECT 69.190 20.580 69.360 20.750 ;
        RECT 69.190 20.220 69.360 20.390 ;
        RECT 69.860 20.755 70.030 20.925 ;
        RECT 69.860 20.395 70.030 20.565 ;
        RECT 71.140 20.755 71.310 20.925 ;
        RECT 71.140 20.395 71.310 20.565 ;
        RECT 72.420 20.755 72.590 20.925 ;
        RECT 72.420 20.395 72.590 20.565 ;
        RECT 74.700 20.755 74.870 20.925 ;
        RECT 74.700 20.395 74.870 20.565 ;
        RECT 76.980 20.755 77.150 20.925 ;
        RECT 76.980 20.395 77.150 20.565 ;
        RECT 78.260 20.755 78.430 20.925 ;
        RECT 78.260 20.395 78.430 20.565 ;
        RECT 79.540 20.755 79.710 20.925 ;
        RECT 79.540 20.395 79.710 20.565 ;
        RECT 80.820 20.755 80.990 20.925 ;
        RECT 80.820 20.395 80.990 20.565 ;
        RECT 82.100 20.755 82.270 20.925 ;
        RECT 82.100 20.395 82.270 20.565 ;
        RECT 84.380 20.755 84.550 20.925 ;
        RECT 84.380 20.395 84.550 20.565 ;
        RECT 86.660 20.755 86.830 20.925 ;
        RECT 86.660 20.395 86.830 20.565 ;
        RECT 87.940 20.755 88.110 20.925 ;
        RECT 87.940 20.395 88.110 20.565 ;
        RECT 89.220 20.755 89.390 20.925 ;
        RECT 89.220 20.395 89.390 20.565 ;
        RECT 135.120 21.840 135.290 22.010 ;
        RECT 144.200 21.840 144.370 22.010 ;
        RECT 135.120 21.480 135.290 21.650 ;
        RECT 89.890 20.940 90.060 21.110 ;
        RECT 89.890 20.580 90.060 20.750 ;
        RECT 89.890 20.220 90.060 20.390 ;
        RECT 69.190 19.860 69.360 20.030 ;
        RECT 69.190 19.500 69.360 19.670 ;
        RECT 70.245 19.740 70.415 19.910 ;
        RECT 70.605 19.740 70.775 19.910 ;
        RECT 70.965 19.740 71.135 19.910 ;
        RECT 71.325 19.740 71.495 19.910 ;
        RECT 71.685 19.740 71.855 19.910 ;
        RECT 72.045 19.740 72.215 19.910 ;
        RECT 72.840 19.740 73.010 19.910 ;
        RECT 73.200 19.740 73.370 19.910 ;
        RECT 73.560 19.740 73.730 19.910 ;
        RECT 73.920 19.740 74.090 19.910 ;
        RECT 74.280 19.740 74.450 19.910 ;
        RECT 75.120 19.740 75.290 19.910 ;
        RECT 75.480 19.740 75.650 19.910 ;
        RECT 75.840 19.740 76.010 19.910 ;
        RECT 76.200 19.740 76.370 19.910 ;
        RECT 76.560 19.740 76.730 19.910 ;
        RECT 77.365 19.740 77.535 19.910 ;
        RECT 77.725 19.740 77.895 19.910 ;
        RECT 78.085 19.740 78.255 19.910 ;
        RECT 78.445 19.740 78.615 19.910 ;
        RECT 78.805 19.740 78.975 19.910 ;
        RECT 79.165 19.740 79.335 19.910 ;
        RECT 79.925 19.740 80.095 19.910 ;
        RECT 80.285 19.740 80.455 19.910 ;
        RECT 80.645 19.740 80.815 19.910 ;
        RECT 81.005 19.740 81.175 19.910 ;
        RECT 81.365 19.740 81.535 19.910 ;
        RECT 81.725 19.740 81.895 19.910 ;
        RECT 87.045 19.740 87.215 19.910 ;
        RECT 87.405 19.740 87.575 19.910 ;
        RECT 87.765 19.740 87.935 19.910 ;
        RECT 88.125 19.740 88.295 19.910 ;
        RECT 88.485 19.740 88.655 19.910 ;
        RECT 88.845 19.740 89.015 19.910 ;
        RECT 89.890 19.860 90.060 20.030 ;
        RECT 89.890 19.500 90.060 19.670 ;
        RECT 69.540 19.190 69.710 19.360 ;
        RECT 69.900 19.190 70.070 19.360 ;
        RECT 70.260 19.190 70.430 19.360 ;
        RECT 70.620 19.190 70.790 19.360 ;
        RECT 70.980 19.190 71.150 19.360 ;
        RECT 71.340 19.190 71.510 19.360 ;
        RECT 71.700 19.190 71.870 19.360 ;
        RECT 72.060 19.190 72.230 19.360 ;
        RECT 72.420 19.190 72.590 19.360 ;
        RECT 72.780 19.190 72.950 19.360 ;
        RECT 73.140 19.190 73.310 19.360 ;
        RECT 73.500 19.190 73.670 19.360 ;
        RECT 73.860 19.190 74.030 19.360 ;
        RECT 74.220 19.190 74.390 19.360 ;
        RECT 74.580 19.190 74.750 19.360 ;
        RECT 74.940 19.190 75.110 19.360 ;
        RECT 75.300 19.190 75.470 19.360 ;
        RECT 75.660 19.190 75.830 19.360 ;
        RECT 76.020 19.190 76.190 19.360 ;
        RECT 76.380 19.190 76.550 19.360 ;
        RECT 76.740 19.190 76.910 19.360 ;
        RECT 77.100 19.190 77.270 19.360 ;
        RECT 77.460 19.190 77.630 19.360 ;
        RECT 77.820 19.190 77.990 19.360 ;
        RECT 78.180 19.190 78.350 19.360 ;
        RECT 78.540 19.190 78.710 19.360 ;
        RECT 78.900 19.190 79.070 19.360 ;
        RECT 79.260 19.190 79.430 19.360 ;
        RECT 79.620 19.190 79.790 19.360 ;
        RECT 79.980 19.190 80.150 19.360 ;
        RECT 80.340 19.190 80.510 19.360 ;
        RECT 80.700 19.190 80.870 19.360 ;
        RECT 81.060 19.190 81.230 19.360 ;
        RECT 81.420 19.190 81.590 19.360 ;
        RECT 81.780 19.190 81.950 19.360 ;
        RECT 82.140 19.190 82.310 19.360 ;
        RECT 82.500 19.190 82.670 19.360 ;
        RECT 82.860 19.190 83.030 19.360 ;
        RECT 83.220 19.190 83.390 19.360 ;
        RECT 83.580 19.190 83.750 19.360 ;
        RECT 83.940 19.190 84.110 19.360 ;
        RECT 84.300 19.190 84.470 19.360 ;
        RECT 84.660 19.190 84.830 19.360 ;
        RECT 85.020 19.190 85.190 19.360 ;
        RECT 85.380 19.190 85.550 19.360 ;
        RECT 85.740 19.190 85.910 19.360 ;
        RECT 86.100 19.190 86.270 19.360 ;
        RECT 86.460 19.190 86.630 19.360 ;
        RECT 86.820 19.190 86.990 19.360 ;
        RECT 87.180 19.190 87.350 19.360 ;
        RECT 87.540 19.190 87.710 19.360 ;
        RECT 87.900 19.190 88.070 19.360 ;
        RECT 88.260 19.190 88.430 19.360 ;
        RECT 88.620 19.190 88.790 19.360 ;
        RECT 88.980 19.190 89.150 19.360 ;
        RECT 89.340 19.190 89.510 19.360 ;
        RECT 94.490 21.075 94.660 21.245 ;
        RECT 94.850 21.075 95.020 21.245 ;
        RECT 95.210 21.075 95.380 21.245 ;
        RECT 95.570 21.075 95.740 21.245 ;
        RECT 95.930 21.075 96.100 21.245 ;
        RECT 96.290 21.075 96.460 21.245 ;
        RECT 96.650 21.075 96.820 21.245 ;
        RECT 97.010 21.075 97.180 21.245 ;
        RECT 97.370 21.075 97.540 21.245 ;
        RECT 97.730 21.075 97.900 21.245 ;
        RECT 98.090 21.075 98.260 21.245 ;
        RECT 98.450 21.075 98.620 21.245 ;
        RECT 98.810 21.075 98.980 21.245 ;
        RECT 99.170 21.075 99.340 21.245 ;
        RECT 99.530 21.075 99.700 21.245 ;
        RECT 99.890 21.075 100.060 21.245 ;
        RECT 100.250 21.075 100.420 21.245 ;
        RECT 100.610 21.075 100.780 21.245 ;
        RECT 100.970 21.075 101.140 21.245 ;
        RECT 101.330 21.075 101.500 21.245 ;
        RECT 101.690 21.075 101.860 21.245 ;
        RECT 102.050 21.075 102.220 21.245 ;
        RECT 102.410 21.075 102.580 21.245 ;
        RECT 102.770 21.075 102.940 21.245 ;
        RECT 103.130 21.075 103.300 21.245 ;
        RECT 103.490 21.075 103.660 21.245 ;
        RECT 103.850 21.075 104.020 21.245 ;
        RECT 104.210 21.075 104.380 21.245 ;
        RECT 104.570 21.075 104.740 21.245 ;
        RECT 104.930 21.075 105.100 21.245 ;
        RECT 105.290 21.075 105.460 21.245 ;
        RECT 105.650 21.075 105.820 21.245 ;
        RECT 106.010 21.075 106.180 21.245 ;
        RECT 106.370 21.075 106.540 21.245 ;
        RECT 106.730 21.075 106.900 21.245 ;
        RECT 107.090 21.075 107.260 21.245 ;
        RECT 107.450 21.075 107.620 21.245 ;
        RECT 107.810 21.075 107.980 21.245 ;
        RECT 108.170 21.075 108.340 21.245 ;
        RECT 108.530 21.075 108.700 21.245 ;
        RECT 108.890 21.075 109.060 21.245 ;
        RECT 109.250 21.075 109.420 21.245 ;
        RECT 109.610 21.075 109.780 21.245 ;
        RECT 109.970 21.075 110.140 21.245 ;
        RECT 110.330 21.075 110.500 21.245 ;
        RECT 110.690 21.075 110.860 21.245 ;
        RECT 111.050 21.075 111.220 21.245 ;
        RECT 111.410 21.075 111.580 21.245 ;
        RECT 111.770 21.075 111.940 21.245 ;
        RECT 112.130 21.075 112.300 21.245 ;
        RECT 112.490 21.075 112.660 21.245 ;
        RECT 112.850 21.075 113.020 21.245 ;
        RECT 113.210 21.075 113.380 21.245 ;
        RECT 113.570 21.075 113.740 21.245 ;
        RECT 113.930 21.075 114.100 21.245 ;
        RECT 114.290 21.075 114.460 21.245 ;
        RECT 114.650 21.075 114.820 21.245 ;
        RECT 115.010 21.075 115.180 21.245 ;
        RECT 115.370 21.075 115.540 21.245 ;
        RECT 115.730 21.075 115.900 21.245 ;
        RECT 116.090 21.075 116.260 21.245 ;
        RECT 116.450 21.075 116.620 21.245 ;
        RECT 116.810 21.075 116.980 21.245 ;
        RECT 117.170 21.075 117.340 21.245 ;
        RECT 117.530 21.075 117.700 21.245 ;
        RECT 117.890 21.075 118.060 21.245 ;
        RECT 94.140 20.775 94.310 20.945 ;
        RECT 118.280 20.775 118.450 20.945 ;
        RECT 94.140 20.415 94.310 20.585 ;
        RECT 94.140 20.055 94.310 20.225 ;
        RECT 94.810 20.280 94.980 20.450 ;
        RECT 97.090 20.280 97.260 20.450 ;
        RECT 99.370 20.280 99.540 20.450 ;
        RECT 101.650 20.280 101.820 20.450 ;
        RECT 103.930 20.280 104.100 20.450 ;
        RECT 106.210 20.280 106.380 20.450 ;
        RECT 108.490 20.280 108.660 20.450 ;
        RECT 110.770 20.280 110.940 20.450 ;
        RECT 113.050 20.280 113.220 20.450 ;
        RECT 115.330 20.280 115.500 20.450 ;
        RECT 117.610 20.280 117.780 20.450 ;
        RECT 118.280 20.415 118.450 20.585 ;
        RECT 118.280 20.055 118.450 20.225 ;
        RECT 94.140 19.695 94.310 19.865 ;
        RECT 95.230 19.695 95.400 19.865 ;
        RECT 95.590 19.695 95.760 19.865 ;
        RECT 95.950 19.695 96.120 19.865 ;
        RECT 96.310 19.695 96.480 19.865 ;
        RECT 96.670 19.695 96.840 19.865 ;
        RECT 97.510 19.695 97.680 19.865 ;
        RECT 97.870 19.695 98.040 19.865 ;
        RECT 98.230 19.695 98.400 19.865 ;
        RECT 98.590 19.695 98.760 19.865 ;
        RECT 98.950 19.695 99.120 19.865 ;
        RECT 99.790 19.695 99.960 19.865 ;
        RECT 100.150 19.695 100.320 19.865 ;
        RECT 100.510 19.695 100.680 19.865 ;
        RECT 100.870 19.695 101.040 19.865 ;
        RECT 101.230 19.695 101.400 19.865 ;
        RECT 102.070 19.695 102.240 19.865 ;
        RECT 102.430 19.695 102.600 19.865 ;
        RECT 102.790 19.695 102.960 19.865 ;
        RECT 103.150 19.695 103.320 19.865 ;
        RECT 103.510 19.695 103.680 19.865 ;
        RECT 104.350 19.695 104.520 19.865 ;
        RECT 104.710 19.695 104.880 19.865 ;
        RECT 105.070 19.695 105.240 19.865 ;
        RECT 105.430 19.695 105.600 19.865 ;
        RECT 105.790 19.695 105.960 19.865 ;
        RECT 106.630 19.695 106.800 19.865 ;
        RECT 106.990 19.695 107.160 19.865 ;
        RECT 107.350 19.695 107.520 19.865 ;
        RECT 107.710 19.695 107.880 19.865 ;
        RECT 108.070 19.695 108.240 19.865 ;
        RECT 108.910 19.695 109.080 19.865 ;
        RECT 109.270 19.695 109.440 19.865 ;
        RECT 109.630 19.695 109.800 19.865 ;
        RECT 109.990 19.695 110.160 19.865 ;
        RECT 110.350 19.695 110.520 19.865 ;
        RECT 111.190 19.695 111.360 19.865 ;
        RECT 111.550 19.695 111.720 19.865 ;
        RECT 111.910 19.695 112.080 19.865 ;
        RECT 112.270 19.695 112.440 19.865 ;
        RECT 112.630 19.695 112.800 19.865 ;
        RECT 113.470 19.695 113.640 19.865 ;
        RECT 113.830 19.695 114.000 19.865 ;
        RECT 114.190 19.695 114.360 19.865 ;
        RECT 114.550 19.695 114.720 19.865 ;
        RECT 114.910 19.695 115.080 19.865 ;
        RECT 115.750 19.695 115.920 19.865 ;
        RECT 116.110 19.695 116.280 19.865 ;
        RECT 116.470 19.695 116.640 19.865 ;
        RECT 116.830 19.695 117.000 19.865 ;
        RECT 117.190 19.695 117.360 19.865 ;
        RECT 118.280 19.695 118.450 19.865 ;
        RECT 94.140 19.335 94.310 19.505 ;
        RECT 94.140 18.975 94.310 19.145 ;
        RECT 118.280 19.335 118.450 19.505 ;
        RECT 118.280 18.975 118.450 19.145 ;
        RECT 135.120 21.120 135.290 21.290 ;
        RECT 135.120 20.760 135.290 20.930 ;
        RECT 135.120 20.400 135.290 20.570 ;
        RECT 135.120 20.040 135.290 20.210 ;
        RECT 135.120 19.680 135.290 19.850 ;
        RECT 135.790 21.315 135.960 21.485 ;
        RECT 135.790 20.955 135.960 21.125 ;
        RECT 135.790 20.595 135.960 20.765 ;
        RECT 135.790 20.235 135.960 20.405 ;
        RECT 135.790 19.875 135.960 20.045 ;
        RECT 136.220 21.315 136.390 21.485 ;
        RECT 136.220 20.955 136.390 21.125 ;
        RECT 136.220 20.595 136.390 20.765 ;
        RECT 136.220 20.235 136.390 20.405 ;
        RECT 136.220 19.875 136.390 20.045 ;
        RECT 136.650 21.315 136.820 21.485 ;
        RECT 136.650 20.955 136.820 21.125 ;
        RECT 136.650 20.595 136.820 20.765 ;
        RECT 136.650 20.235 136.820 20.405 ;
        RECT 136.650 19.875 136.820 20.045 ;
        RECT 137.080 21.315 137.250 21.485 ;
        RECT 137.080 20.955 137.250 21.125 ;
        RECT 137.080 20.595 137.250 20.765 ;
        RECT 137.080 20.235 137.250 20.405 ;
        RECT 137.080 19.875 137.250 20.045 ;
        RECT 137.510 21.315 137.680 21.485 ;
        RECT 137.510 20.955 137.680 21.125 ;
        RECT 137.510 20.595 137.680 20.765 ;
        RECT 137.510 20.235 137.680 20.405 ;
        RECT 137.510 19.875 137.680 20.045 ;
        RECT 137.940 21.315 138.110 21.485 ;
        RECT 137.940 20.955 138.110 21.125 ;
        RECT 137.940 20.595 138.110 20.765 ;
        RECT 137.940 20.235 138.110 20.405 ;
        RECT 137.940 19.875 138.110 20.045 ;
        RECT 138.370 21.315 138.540 21.485 ;
        RECT 138.370 20.955 138.540 21.125 ;
        RECT 138.370 20.595 138.540 20.765 ;
        RECT 138.370 20.235 138.540 20.405 ;
        RECT 138.370 19.875 138.540 20.045 ;
        RECT 138.800 21.315 138.970 21.485 ;
        RECT 138.800 20.955 138.970 21.125 ;
        RECT 138.800 20.595 138.970 20.765 ;
        RECT 138.800 20.235 138.970 20.405 ;
        RECT 138.800 19.875 138.970 20.045 ;
        RECT 139.230 21.315 139.400 21.485 ;
        RECT 139.230 20.955 139.400 21.125 ;
        RECT 139.230 20.595 139.400 20.765 ;
        RECT 139.230 20.235 139.400 20.405 ;
        RECT 139.230 19.875 139.400 20.045 ;
        RECT 139.660 21.315 139.830 21.485 ;
        RECT 139.660 20.955 139.830 21.125 ;
        RECT 139.660 20.595 139.830 20.765 ;
        RECT 139.660 20.235 139.830 20.405 ;
        RECT 139.660 19.875 139.830 20.045 ;
        RECT 140.090 21.315 140.260 21.485 ;
        RECT 140.090 20.955 140.260 21.125 ;
        RECT 140.090 20.595 140.260 20.765 ;
        RECT 140.090 20.235 140.260 20.405 ;
        RECT 140.090 19.875 140.260 20.045 ;
        RECT 140.520 21.315 140.690 21.485 ;
        RECT 140.520 20.955 140.690 21.125 ;
        RECT 140.520 20.595 140.690 20.765 ;
        RECT 140.520 20.235 140.690 20.405 ;
        RECT 140.520 19.875 140.690 20.045 ;
        RECT 140.950 21.315 141.120 21.485 ;
        RECT 140.950 20.955 141.120 21.125 ;
        RECT 140.950 20.595 141.120 20.765 ;
        RECT 140.950 20.235 141.120 20.405 ;
        RECT 140.950 19.875 141.120 20.045 ;
        RECT 141.380 21.315 141.550 21.485 ;
        RECT 141.380 20.955 141.550 21.125 ;
        RECT 141.380 20.595 141.550 20.765 ;
        RECT 141.380 20.235 141.550 20.405 ;
        RECT 141.380 19.875 141.550 20.045 ;
        RECT 141.810 21.315 141.980 21.485 ;
        RECT 141.810 20.955 141.980 21.125 ;
        RECT 141.810 20.595 141.980 20.765 ;
        RECT 141.810 20.235 141.980 20.405 ;
        RECT 141.810 19.875 141.980 20.045 ;
        RECT 142.240 21.315 142.410 21.485 ;
        RECT 142.240 20.955 142.410 21.125 ;
        RECT 142.240 20.595 142.410 20.765 ;
        RECT 142.240 20.235 142.410 20.405 ;
        RECT 142.240 19.875 142.410 20.045 ;
        RECT 142.670 21.315 142.840 21.485 ;
        RECT 142.670 20.955 142.840 21.125 ;
        RECT 142.670 20.595 142.840 20.765 ;
        RECT 142.670 20.235 142.840 20.405 ;
        RECT 142.670 19.875 142.840 20.045 ;
        RECT 143.100 21.315 143.270 21.485 ;
        RECT 143.100 20.955 143.270 21.125 ;
        RECT 143.100 20.595 143.270 20.765 ;
        RECT 143.100 20.235 143.270 20.405 ;
        RECT 143.100 19.875 143.270 20.045 ;
        RECT 143.530 21.315 143.700 21.485 ;
        RECT 143.530 20.955 143.700 21.125 ;
        RECT 143.530 20.595 143.700 20.765 ;
        RECT 143.530 20.235 143.700 20.405 ;
        RECT 143.530 19.875 143.700 20.045 ;
        RECT 144.200 21.480 144.370 21.650 ;
        RECT 144.200 21.120 144.370 21.290 ;
        RECT 144.200 20.760 144.370 20.930 ;
        RECT 144.200 20.400 144.370 20.570 ;
        RECT 144.200 20.040 144.370 20.210 ;
        RECT 144.200 19.680 144.370 19.850 ;
        RECT 135.120 19.320 135.290 19.490 ;
        RECT 136.040 19.260 136.210 19.430 ;
        RECT 136.400 19.260 136.570 19.430 ;
        RECT 136.900 19.260 137.070 19.430 ;
        RECT 137.260 19.260 137.430 19.430 ;
        RECT 137.760 19.260 137.930 19.430 ;
        RECT 138.120 19.260 138.290 19.430 ;
        RECT 138.620 19.260 138.790 19.430 ;
        RECT 138.980 19.260 139.150 19.430 ;
        RECT 139.480 19.260 139.650 19.430 ;
        RECT 139.840 19.260 140.010 19.430 ;
        RECT 140.340 19.260 140.510 19.430 ;
        RECT 140.700 19.260 140.870 19.430 ;
        RECT 141.200 19.260 141.370 19.430 ;
        RECT 141.560 19.260 141.730 19.430 ;
        RECT 142.060 19.260 142.230 19.430 ;
        RECT 142.420 19.260 142.590 19.430 ;
        RECT 142.920 19.260 143.090 19.430 ;
        RECT 143.280 19.260 143.450 19.430 ;
        RECT 144.200 19.320 144.370 19.490 ;
        RECT 56.330 17.705 56.500 17.875 ;
        RECT 56.690 17.705 56.860 17.875 ;
        RECT 57.050 17.705 57.220 17.875 ;
        RECT 57.410 17.705 57.580 17.875 ;
        RECT 57.770 17.705 57.940 17.875 ;
        RECT 58.130 17.705 58.300 17.875 ;
        RECT 58.490 17.705 58.660 17.875 ;
        RECT 58.850 17.705 59.020 17.875 ;
        RECT 59.210 17.705 59.380 17.875 ;
        RECT 59.570 17.705 59.740 17.875 ;
        RECT 59.930 17.705 60.100 17.875 ;
        RECT 60.290 17.705 60.460 17.875 ;
        RECT 60.650 17.705 60.820 17.875 ;
        RECT 61.010 17.705 61.180 17.875 ;
        RECT 61.370 17.705 61.540 17.875 ;
        RECT 61.730 17.705 61.900 17.875 ;
        RECT 62.090 17.705 62.260 17.875 ;
        RECT 62.450 17.705 62.620 17.875 ;
        RECT 62.810 17.705 62.980 17.875 ;
        RECT 63.170 17.705 63.340 17.875 ;
        RECT 63.530 17.705 63.700 17.875 ;
        RECT 63.890 17.705 64.060 17.875 ;
        RECT 64.250 17.705 64.420 17.875 ;
        RECT 64.610 17.705 64.780 17.875 ;
        RECT 55.980 17.405 56.150 17.575 ;
        RECT 65.000 17.405 65.170 17.575 ;
        RECT 55.980 17.045 56.150 17.215 ;
        RECT 57.070 17.155 57.240 17.325 ;
        RECT 57.430 17.155 57.600 17.325 ;
        RECT 57.790 17.155 57.960 17.325 ;
        RECT 63.190 17.155 63.360 17.325 ;
        RECT 63.550 17.155 63.720 17.325 ;
        RECT 63.910 17.155 64.080 17.325 ;
        RECT 65.000 17.045 65.170 17.215 ;
        RECT 55.980 16.685 56.150 16.855 ;
        RECT 55.980 16.325 56.150 16.495 ;
        RECT 56.650 16.570 56.820 16.740 ;
        RECT 57.430 16.570 57.600 16.740 ;
        RECT 58.210 16.570 58.380 16.740 ;
        RECT 60.490 16.570 60.660 16.740 ;
        RECT 62.770 16.570 62.940 16.740 ;
        RECT 63.550 16.570 63.720 16.740 ;
        RECT 64.330 16.570 64.500 16.740 ;
        RECT 65.000 16.685 65.170 16.855 ;
        RECT 65.000 16.325 65.170 16.495 ;
        RECT 55.980 15.965 56.150 16.135 ;
        RECT 58.630 15.985 58.800 16.155 ;
        RECT 58.990 15.985 59.160 16.155 ;
        RECT 59.350 15.985 59.520 16.155 ;
        RECT 59.710 15.985 59.880 16.155 ;
        RECT 60.070 15.985 60.240 16.155 ;
        RECT 60.910 15.985 61.080 16.155 ;
        RECT 61.270 15.985 61.440 16.155 ;
        RECT 61.630 15.985 61.800 16.155 ;
        RECT 61.990 15.985 62.160 16.155 ;
        RECT 62.350 15.985 62.520 16.155 ;
        RECT 65.000 15.965 65.170 16.135 ;
        RECT 56.330 15.435 56.500 15.605 ;
        RECT 56.690 15.435 56.860 15.605 ;
        RECT 57.050 15.435 57.220 15.605 ;
        RECT 57.410 15.435 57.580 15.605 ;
        RECT 57.770 15.435 57.940 15.605 ;
        RECT 58.130 15.435 58.300 15.605 ;
        RECT 58.490 15.435 58.660 15.605 ;
        RECT 58.850 15.435 59.020 15.605 ;
        RECT 59.210 15.435 59.380 15.605 ;
        RECT 59.570 15.435 59.740 15.605 ;
        RECT 59.930 15.435 60.100 15.605 ;
        RECT 60.290 15.435 60.460 15.605 ;
        RECT 60.650 15.435 60.820 15.605 ;
        RECT 61.010 15.435 61.180 15.605 ;
        RECT 61.370 15.435 61.540 15.605 ;
        RECT 61.730 15.435 61.900 15.605 ;
        RECT 62.090 15.435 62.260 15.605 ;
        RECT 62.450 15.435 62.620 15.605 ;
        RECT 62.810 15.435 62.980 15.605 ;
        RECT 63.170 15.435 63.340 15.605 ;
        RECT 63.530 15.435 63.700 15.605 ;
        RECT 63.890 15.435 64.060 15.605 ;
        RECT 64.250 15.435 64.420 15.605 ;
        RECT 64.610 15.435 64.780 15.605 ;
        RECT 69.540 17.705 69.710 17.875 ;
        RECT 69.900 17.705 70.070 17.875 ;
        RECT 70.260 17.705 70.430 17.875 ;
        RECT 70.620 17.705 70.790 17.875 ;
        RECT 70.980 17.705 71.150 17.875 ;
        RECT 71.340 17.705 71.510 17.875 ;
        RECT 71.700 17.705 71.870 17.875 ;
        RECT 72.060 17.705 72.230 17.875 ;
        RECT 72.420 17.705 72.590 17.875 ;
        RECT 72.780 17.705 72.950 17.875 ;
        RECT 73.140 17.705 73.310 17.875 ;
        RECT 73.500 17.705 73.670 17.875 ;
        RECT 73.860 17.705 74.030 17.875 ;
        RECT 74.220 17.705 74.390 17.875 ;
        RECT 74.580 17.705 74.750 17.875 ;
        RECT 74.940 17.705 75.110 17.875 ;
        RECT 75.300 17.705 75.470 17.875 ;
        RECT 75.660 17.705 75.830 17.875 ;
        RECT 76.020 17.705 76.190 17.875 ;
        RECT 76.380 17.705 76.550 17.875 ;
        RECT 76.740 17.705 76.910 17.875 ;
        RECT 77.100 17.705 77.270 17.875 ;
        RECT 77.460 17.705 77.630 17.875 ;
        RECT 77.820 17.705 77.990 17.875 ;
        RECT 78.180 17.705 78.350 17.875 ;
        RECT 78.540 17.705 78.710 17.875 ;
        RECT 78.900 17.705 79.070 17.875 ;
        RECT 79.260 17.705 79.430 17.875 ;
        RECT 79.620 17.705 79.790 17.875 ;
        RECT 79.980 17.705 80.150 17.875 ;
        RECT 80.340 17.705 80.510 17.875 ;
        RECT 80.700 17.705 80.870 17.875 ;
        RECT 81.060 17.705 81.230 17.875 ;
        RECT 81.420 17.705 81.590 17.875 ;
        RECT 81.780 17.705 81.950 17.875 ;
        RECT 82.140 17.705 82.310 17.875 ;
        RECT 82.500 17.705 82.670 17.875 ;
        RECT 82.860 17.705 83.030 17.875 ;
        RECT 83.220 17.705 83.390 17.875 ;
        RECT 83.580 17.705 83.750 17.875 ;
        RECT 83.940 17.705 84.110 17.875 ;
        RECT 84.300 17.705 84.470 17.875 ;
        RECT 84.660 17.705 84.830 17.875 ;
        RECT 85.020 17.705 85.190 17.875 ;
        RECT 85.380 17.705 85.550 17.875 ;
        RECT 85.740 17.705 85.910 17.875 ;
        RECT 86.100 17.705 86.270 17.875 ;
        RECT 86.460 17.705 86.630 17.875 ;
        RECT 86.820 17.705 86.990 17.875 ;
        RECT 87.180 17.705 87.350 17.875 ;
        RECT 87.540 17.705 87.710 17.875 ;
        RECT 87.900 17.705 88.070 17.875 ;
        RECT 88.260 17.705 88.430 17.875 ;
        RECT 88.620 17.705 88.790 17.875 ;
        RECT 88.980 17.705 89.150 17.875 ;
        RECT 89.340 17.705 89.510 17.875 ;
        RECT 69.190 17.405 69.360 17.575 ;
        RECT 89.890 17.405 90.060 17.575 ;
        RECT 69.190 17.045 69.360 17.215 ;
        RECT 70.245 17.155 70.415 17.325 ;
        RECT 70.605 17.155 70.775 17.325 ;
        RECT 70.965 17.155 71.135 17.325 ;
        RECT 71.325 17.155 71.495 17.325 ;
        RECT 71.685 17.155 71.855 17.325 ;
        RECT 72.045 17.155 72.215 17.325 ;
        RECT 72.840 17.155 73.010 17.325 ;
        RECT 73.200 17.155 73.370 17.325 ;
        RECT 73.560 17.155 73.730 17.325 ;
        RECT 73.920 17.155 74.090 17.325 ;
        RECT 74.280 17.155 74.450 17.325 ;
        RECT 75.120 17.155 75.290 17.325 ;
        RECT 75.480 17.155 75.650 17.325 ;
        RECT 75.840 17.155 76.010 17.325 ;
        RECT 76.200 17.155 76.370 17.325 ;
        RECT 76.560 17.155 76.730 17.325 ;
        RECT 77.365 17.155 77.535 17.325 ;
        RECT 77.725 17.155 77.895 17.325 ;
        RECT 78.085 17.155 78.255 17.325 ;
        RECT 78.445 17.155 78.615 17.325 ;
        RECT 78.805 17.155 78.975 17.325 ;
        RECT 79.165 17.155 79.335 17.325 ;
        RECT 79.925 17.155 80.095 17.325 ;
        RECT 80.285 17.155 80.455 17.325 ;
        RECT 80.645 17.155 80.815 17.325 ;
        RECT 81.005 17.155 81.175 17.325 ;
        RECT 81.365 17.155 81.535 17.325 ;
        RECT 81.725 17.155 81.895 17.325 ;
        RECT 87.045 17.155 87.215 17.325 ;
        RECT 87.405 17.155 87.575 17.325 ;
        RECT 87.765 17.155 87.935 17.325 ;
        RECT 88.125 17.155 88.295 17.325 ;
        RECT 88.485 17.155 88.655 17.325 ;
        RECT 88.845 17.155 89.015 17.325 ;
        RECT 89.890 17.045 90.060 17.215 ;
        RECT 69.190 16.685 69.360 16.855 ;
        RECT 69.190 16.325 69.360 16.495 ;
        RECT 69.860 16.570 70.030 16.740 ;
        RECT 71.140 16.570 71.310 16.740 ;
        RECT 72.420 16.570 72.590 16.740 ;
        RECT 74.700 16.570 74.870 16.740 ;
        RECT 76.980 16.570 77.150 16.740 ;
        RECT 78.260 16.570 78.430 16.740 ;
        RECT 79.540 16.570 79.710 16.740 ;
        RECT 80.820 16.570 80.990 16.740 ;
        RECT 82.100 16.570 82.270 16.740 ;
        RECT 84.380 16.570 84.550 16.740 ;
        RECT 86.660 16.570 86.830 16.740 ;
        RECT 87.940 16.570 88.110 16.740 ;
        RECT 89.220 16.570 89.390 16.740 ;
        RECT 89.890 16.685 90.060 16.855 ;
        RECT 89.890 16.325 90.060 16.495 ;
        RECT 69.190 15.965 69.360 16.135 ;
        RECT 70.245 15.985 70.415 16.155 ;
        RECT 70.605 15.985 70.775 16.155 ;
        RECT 70.965 15.985 71.135 16.155 ;
        RECT 71.325 15.985 71.495 16.155 ;
        RECT 71.685 15.985 71.855 16.155 ;
        RECT 72.045 15.985 72.215 16.155 ;
        RECT 72.840 15.985 73.010 16.155 ;
        RECT 73.200 15.985 73.370 16.155 ;
        RECT 73.560 15.985 73.730 16.155 ;
        RECT 73.920 15.985 74.090 16.155 ;
        RECT 74.280 15.985 74.450 16.155 ;
        RECT 75.120 15.985 75.290 16.155 ;
        RECT 75.480 15.985 75.650 16.155 ;
        RECT 75.840 15.985 76.010 16.155 ;
        RECT 76.200 15.985 76.370 16.155 ;
        RECT 76.560 15.985 76.730 16.155 ;
        RECT 77.365 15.985 77.535 16.155 ;
        RECT 77.725 15.985 77.895 16.155 ;
        RECT 78.085 15.985 78.255 16.155 ;
        RECT 78.445 15.985 78.615 16.155 ;
        RECT 78.805 15.985 78.975 16.155 ;
        RECT 79.165 15.985 79.335 16.155 ;
        RECT 79.925 15.985 80.095 16.155 ;
        RECT 80.285 15.985 80.455 16.155 ;
        RECT 80.645 15.985 80.815 16.155 ;
        RECT 81.005 15.985 81.175 16.155 ;
        RECT 81.365 15.985 81.535 16.155 ;
        RECT 81.725 15.985 81.895 16.155 ;
        RECT 82.520 15.985 82.690 16.155 ;
        RECT 82.880 15.985 83.050 16.155 ;
        RECT 83.240 15.985 83.410 16.155 ;
        RECT 83.600 15.985 83.770 16.155 ;
        RECT 83.960 15.985 84.130 16.155 ;
        RECT 84.800 15.985 84.970 16.155 ;
        RECT 85.160 15.985 85.330 16.155 ;
        RECT 85.520 15.985 85.690 16.155 ;
        RECT 85.880 15.985 86.050 16.155 ;
        RECT 86.240 15.985 86.410 16.155 ;
        RECT 87.045 15.985 87.215 16.155 ;
        RECT 87.405 15.985 87.575 16.155 ;
        RECT 87.765 15.985 87.935 16.155 ;
        RECT 88.125 15.985 88.295 16.155 ;
        RECT 88.485 15.985 88.655 16.155 ;
        RECT 88.845 15.985 89.015 16.155 ;
        RECT 89.890 15.965 90.060 16.135 ;
        RECT 69.540 15.435 69.710 15.605 ;
        RECT 69.900 15.435 70.070 15.605 ;
        RECT 70.260 15.435 70.430 15.605 ;
        RECT 70.620 15.435 70.790 15.605 ;
        RECT 70.980 15.435 71.150 15.605 ;
        RECT 71.340 15.435 71.510 15.605 ;
        RECT 71.700 15.435 71.870 15.605 ;
        RECT 72.060 15.435 72.230 15.605 ;
        RECT 72.420 15.435 72.590 15.605 ;
        RECT 72.780 15.435 72.950 15.605 ;
        RECT 73.140 15.435 73.310 15.605 ;
        RECT 73.500 15.435 73.670 15.605 ;
        RECT 73.860 15.435 74.030 15.605 ;
        RECT 74.220 15.435 74.390 15.605 ;
        RECT 74.580 15.435 74.750 15.605 ;
        RECT 74.940 15.435 75.110 15.605 ;
        RECT 75.300 15.435 75.470 15.605 ;
        RECT 75.660 15.435 75.830 15.605 ;
        RECT 76.020 15.435 76.190 15.605 ;
        RECT 76.380 15.435 76.550 15.605 ;
        RECT 76.740 15.435 76.910 15.605 ;
        RECT 77.100 15.435 77.270 15.605 ;
        RECT 77.460 15.435 77.630 15.605 ;
        RECT 77.820 15.435 77.990 15.605 ;
        RECT 78.180 15.435 78.350 15.605 ;
        RECT 78.540 15.435 78.710 15.605 ;
        RECT 78.900 15.435 79.070 15.605 ;
        RECT 79.260 15.435 79.430 15.605 ;
        RECT 79.620 15.435 79.790 15.605 ;
        RECT 79.980 15.435 80.150 15.605 ;
        RECT 80.340 15.435 80.510 15.605 ;
        RECT 80.700 15.435 80.870 15.605 ;
        RECT 81.060 15.435 81.230 15.605 ;
        RECT 81.420 15.435 81.590 15.605 ;
        RECT 81.780 15.435 81.950 15.605 ;
        RECT 82.140 15.435 82.310 15.605 ;
        RECT 82.500 15.435 82.670 15.605 ;
        RECT 82.860 15.435 83.030 15.605 ;
        RECT 83.220 15.435 83.390 15.605 ;
        RECT 83.580 15.435 83.750 15.605 ;
        RECT 83.940 15.435 84.110 15.605 ;
        RECT 84.300 15.435 84.470 15.605 ;
        RECT 84.660 15.435 84.830 15.605 ;
        RECT 85.020 15.435 85.190 15.605 ;
        RECT 85.380 15.435 85.550 15.605 ;
        RECT 85.740 15.435 85.910 15.605 ;
        RECT 86.100 15.435 86.270 15.605 ;
        RECT 86.460 15.435 86.630 15.605 ;
        RECT 86.820 15.435 86.990 15.605 ;
        RECT 87.180 15.435 87.350 15.605 ;
        RECT 87.540 15.435 87.710 15.605 ;
        RECT 87.900 15.435 88.070 15.605 ;
        RECT 88.260 15.435 88.430 15.605 ;
        RECT 88.620 15.435 88.790 15.605 ;
        RECT 88.980 15.435 89.150 15.605 ;
        RECT 89.340 15.435 89.510 15.605 ;
        RECT 94.140 17.505 94.310 17.675 ;
        RECT 94.140 17.145 94.310 17.315 ;
        RECT 94.140 16.785 94.310 16.955 ;
        RECT 118.280 17.505 118.450 17.675 ;
        RECT 118.280 17.145 118.450 17.315 ;
        RECT 94.140 16.425 94.310 16.595 ;
        RECT 95.230 16.565 95.400 16.735 ;
        RECT 95.590 16.565 95.760 16.735 ;
        RECT 95.950 16.565 96.120 16.735 ;
        RECT 96.310 16.565 96.480 16.735 ;
        RECT 96.670 16.565 96.840 16.735 ;
        RECT 97.510 16.565 97.680 16.735 ;
        RECT 97.870 16.565 98.040 16.735 ;
        RECT 98.230 16.565 98.400 16.735 ;
        RECT 98.590 16.565 98.760 16.735 ;
        RECT 98.950 16.565 99.120 16.735 ;
        RECT 99.790 16.565 99.960 16.735 ;
        RECT 100.150 16.565 100.320 16.735 ;
        RECT 100.510 16.565 100.680 16.735 ;
        RECT 100.870 16.565 101.040 16.735 ;
        RECT 101.230 16.565 101.400 16.735 ;
        RECT 102.070 16.565 102.240 16.735 ;
        RECT 102.430 16.565 102.600 16.735 ;
        RECT 102.790 16.565 102.960 16.735 ;
        RECT 103.150 16.565 103.320 16.735 ;
        RECT 103.510 16.565 103.680 16.735 ;
        RECT 104.350 16.565 104.520 16.735 ;
        RECT 104.710 16.565 104.880 16.735 ;
        RECT 105.070 16.565 105.240 16.735 ;
        RECT 105.430 16.565 105.600 16.735 ;
        RECT 105.790 16.565 105.960 16.735 ;
        RECT 106.630 16.565 106.800 16.735 ;
        RECT 106.990 16.565 107.160 16.735 ;
        RECT 107.350 16.565 107.520 16.735 ;
        RECT 107.710 16.565 107.880 16.735 ;
        RECT 108.070 16.565 108.240 16.735 ;
        RECT 108.910 16.565 109.080 16.735 ;
        RECT 109.270 16.565 109.440 16.735 ;
        RECT 109.630 16.565 109.800 16.735 ;
        RECT 109.990 16.565 110.160 16.735 ;
        RECT 110.350 16.565 110.520 16.735 ;
        RECT 111.190 16.565 111.360 16.735 ;
        RECT 111.550 16.565 111.720 16.735 ;
        RECT 111.910 16.565 112.080 16.735 ;
        RECT 112.270 16.565 112.440 16.735 ;
        RECT 112.630 16.565 112.800 16.735 ;
        RECT 113.470 16.565 113.640 16.735 ;
        RECT 113.830 16.565 114.000 16.735 ;
        RECT 114.190 16.565 114.360 16.735 ;
        RECT 114.550 16.565 114.720 16.735 ;
        RECT 114.910 16.565 115.080 16.735 ;
        RECT 115.750 16.565 115.920 16.735 ;
        RECT 116.110 16.565 116.280 16.735 ;
        RECT 116.470 16.565 116.640 16.735 ;
        RECT 116.830 16.565 117.000 16.735 ;
        RECT 117.190 16.565 117.360 16.735 ;
        RECT 118.280 16.785 118.450 16.955 ;
        RECT 118.280 16.425 118.450 16.595 ;
        RECT 94.140 16.065 94.310 16.235 ;
        RECT 94.140 15.705 94.310 15.875 ;
        RECT 94.140 15.345 94.310 15.515 ;
        RECT 94.810 15.910 94.980 16.080 ;
        RECT 94.810 15.550 94.980 15.720 ;
        RECT 97.090 15.910 97.260 16.080 ;
        RECT 97.090 15.550 97.260 15.720 ;
        RECT 99.370 15.910 99.540 16.080 ;
        RECT 99.370 15.550 99.540 15.720 ;
        RECT 101.650 15.910 101.820 16.080 ;
        RECT 101.650 15.550 101.820 15.720 ;
        RECT 103.930 15.910 104.100 16.080 ;
        RECT 103.930 15.550 104.100 15.720 ;
        RECT 106.210 15.910 106.380 16.080 ;
        RECT 106.210 15.550 106.380 15.720 ;
        RECT 108.490 15.910 108.660 16.080 ;
        RECT 108.490 15.550 108.660 15.720 ;
        RECT 110.770 15.910 110.940 16.080 ;
        RECT 110.770 15.550 110.940 15.720 ;
        RECT 113.050 15.910 113.220 16.080 ;
        RECT 113.050 15.550 113.220 15.720 ;
        RECT 115.330 15.910 115.500 16.080 ;
        RECT 115.330 15.550 115.500 15.720 ;
        RECT 117.610 15.910 117.780 16.080 ;
        RECT 117.610 15.550 117.780 15.720 ;
        RECT 118.280 16.065 118.450 16.235 ;
        RECT 118.280 15.705 118.450 15.875 ;
        RECT 135.120 17.825 135.290 17.995 ;
        RECT 135.120 17.465 135.290 17.635 ;
        RECT 136.040 17.580 136.210 17.750 ;
        RECT 136.400 17.580 136.570 17.750 ;
        RECT 136.900 17.580 137.070 17.750 ;
        RECT 137.260 17.580 137.430 17.750 ;
        RECT 137.760 17.580 137.930 17.750 ;
        RECT 138.120 17.580 138.290 17.750 ;
        RECT 138.620 17.580 138.790 17.750 ;
        RECT 138.980 17.580 139.150 17.750 ;
        RECT 139.480 17.580 139.650 17.750 ;
        RECT 139.840 17.580 140.010 17.750 ;
        RECT 140.340 17.580 140.510 17.750 ;
        RECT 140.700 17.580 140.870 17.750 ;
        RECT 141.200 17.580 141.370 17.750 ;
        RECT 141.560 17.580 141.730 17.750 ;
        RECT 142.060 17.580 142.230 17.750 ;
        RECT 142.420 17.580 142.590 17.750 ;
        RECT 142.920 17.580 143.090 17.750 ;
        RECT 143.280 17.580 143.450 17.750 ;
        RECT 144.200 17.825 144.370 17.995 ;
        RECT 144.200 17.465 144.370 17.635 ;
        RECT 135.120 17.105 135.290 17.275 ;
        RECT 135.120 16.745 135.290 16.915 ;
        RECT 135.120 16.385 135.290 16.555 ;
        RECT 135.790 16.925 135.960 17.095 ;
        RECT 135.790 16.565 135.960 16.735 ;
        RECT 136.220 16.925 136.390 17.095 ;
        RECT 136.220 16.565 136.390 16.735 ;
        RECT 136.650 16.925 136.820 17.095 ;
        RECT 136.650 16.565 136.820 16.735 ;
        RECT 137.080 16.925 137.250 17.095 ;
        RECT 137.080 16.565 137.250 16.735 ;
        RECT 137.510 16.925 137.680 17.095 ;
        RECT 137.510 16.565 137.680 16.735 ;
        RECT 137.940 16.925 138.110 17.095 ;
        RECT 137.940 16.565 138.110 16.735 ;
        RECT 138.370 16.925 138.540 17.095 ;
        RECT 138.370 16.565 138.540 16.735 ;
        RECT 138.800 16.925 138.970 17.095 ;
        RECT 138.800 16.565 138.970 16.735 ;
        RECT 139.230 16.925 139.400 17.095 ;
        RECT 139.230 16.565 139.400 16.735 ;
        RECT 139.660 16.925 139.830 17.095 ;
        RECT 139.660 16.565 139.830 16.735 ;
        RECT 140.090 16.925 140.260 17.095 ;
        RECT 140.090 16.565 140.260 16.735 ;
        RECT 140.520 16.925 140.690 17.095 ;
        RECT 140.520 16.565 140.690 16.735 ;
        RECT 140.950 16.925 141.120 17.095 ;
        RECT 140.950 16.565 141.120 16.735 ;
        RECT 141.380 16.925 141.550 17.095 ;
        RECT 141.380 16.565 141.550 16.735 ;
        RECT 141.810 16.925 141.980 17.095 ;
        RECT 141.810 16.565 141.980 16.735 ;
        RECT 142.240 16.925 142.410 17.095 ;
        RECT 142.240 16.565 142.410 16.735 ;
        RECT 142.670 16.925 142.840 17.095 ;
        RECT 142.670 16.565 142.840 16.735 ;
        RECT 143.100 16.925 143.270 17.095 ;
        RECT 143.100 16.565 143.270 16.735 ;
        RECT 143.530 16.925 143.700 17.095 ;
        RECT 143.530 16.565 143.700 16.735 ;
        RECT 144.200 17.105 144.370 17.275 ;
        RECT 144.200 16.745 144.370 16.915 ;
        RECT 144.200 16.385 144.370 16.555 ;
        RECT 135.120 16.025 135.290 16.195 ;
        RECT 144.200 16.025 144.370 16.195 ;
        RECT 135.470 15.725 135.640 15.895 ;
        RECT 135.830 15.725 136.000 15.895 ;
        RECT 136.190 15.725 136.360 15.895 ;
        RECT 136.550 15.725 136.720 15.895 ;
        RECT 136.910 15.725 137.080 15.895 ;
        RECT 137.270 15.725 137.440 15.895 ;
        RECT 137.630 15.725 137.800 15.895 ;
        RECT 137.990 15.725 138.160 15.895 ;
        RECT 138.350 15.725 138.520 15.895 ;
        RECT 138.710 15.725 138.880 15.895 ;
        RECT 139.070 15.725 139.240 15.895 ;
        RECT 139.430 15.725 139.600 15.895 ;
        RECT 139.790 15.725 139.960 15.895 ;
        RECT 140.150 15.725 140.320 15.895 ;
        RECT 140.510 15.725 140.680 15.895 ;
        RECT 140.870 15.725 141.040 15.895 ;
        RECT 141.230 15.725 141.400 15.895 ;
        RECT 141.590 15.725 141.760 15.895 ;
        RECT 141.950 15.725 142.120 15.895 ;
        RECT 142.310 15.725 142.480 15.895 ;
        RECT 142.670 15.725 142.840 15.895 ;
        RECT 143.030 15.725 143.200 15.895 ;
        RECT 143.390 15.725 143.560 15.895 ;
        RECT 143.750 15.725 143.920 15.895 ;
        RECT 118.280 15.345 118.450 15.515 ;
        RECT 94.140 14.985 94.310 15.155 ;
        RECT 118.280 14.985 118.450 15.155 ;
        RECT 94.490 14.685 94.660 14.855 ;
        RECT 94.850 14.685 95.020 14.855 ;
        RECT 95.210 14.685 95.380 14.855 ;
        RECT 95.570 14.685 95.740 14.855 ;
        RECT 95.930 14.685 96.100 14.855 ;
        RECT 96.290 14.685 96.460 14.855 ;
        RECT 96.650 14.685 96.820 14.855 ;
        RECT 97.010 14.685 97.180 14.855 ;
        RECT 97.370 14.685 97.540 14.855 ;
        RECT 97.730 14.685 97.900 14.855 ;
        RECT 98.090 14.685 98.260 14.855 ;
        RECT 98.450 14.685 98.620 14.855 ;
        RECT 98.810 14.685 98.980 14.855 ;
        RECT 99.170 14.685 99.340 14.855 ;
        RECT 99.530 14.685 99.700 14.855 ;
        RECT 99.890 14.685 100.060 14.855 ;
        RECT 100.250 14.685 100.420 14.855 ;
        RECT 100.610 14.685 100.780 14.855 ;
        RECT 100.970 14.685 101.140 14.855 ;
        RECT 101.330 14.685 101.500 14.855 ;
        RECT 101.690 14.685 101.860 14.855 ;
        RECT 102.050 14.685 102.220 14.855 ;
        RECT 102.410 14.685 102.580 14.855 ;
        RECT 102.770 14.685 102.940 14.855 ;
        RECT 103.130 14.685 103.300 14.855 ;
        RECT 103.490 14.685 103.660 14.855 ;
        RECT 103.850 14.685 104.020 14.855 ;
        RECT 104.210 14.685 104.380 14.855 ;
        RECT 104.570 14.685 104.740 14.855 ;
        RECT 104.930 14.685 105.100 14.855 ;
        RECT 105.290 14.685 105.460 14.855 ;
        RECT 105.650 14.685 105.820 14.855 ;
        RECT 106.010 14.685 106.180 14.855 ;
        RECT 106.370 14.685 106.540 14.855 ;
        RECT 106.730 14.685 106.900 14.855 ;
        RECT 107.090 14.685 107.260 14.855 ;
        RECT 107.450 14.685 107.620 14.855 ;
        RECT 107.810 14.685 107.980 14.855 ;
        RECT 108.170 14.685 108.340 14.855 ;
        RECT 108.530 14.685 108.700 14.855 ;
        RECT 108.890 14.685 109.060 14.855 ;
        RECT 109.250 14.685 109.420 14.855 ;
        RECT 109.610 14.685 109.780 14.855 ;
        RECT 109.970 14.685 110.140 14.855 ;
        RECT 110.330 14.685 110.500 14.855 ;
        RECT 110.690 14.685 110.860 14.855 ;
        RECT 111.050 14.685 111.220 14.855 ;
        RECT 111.410 14.685 111.580 14.855 ;
        RECT 111.770 14.685 111.940 14.855 ;
        RECT 112.130 14.685 112.300 14.855 ;
        RECT 112.490 14.685 112.660 14.855 ;
        RECT 112.850 14.685 113.020 14.855 ;
        RECT 113.210 14.685 113.380 14.855 ;
        RECT 113.570 14.685 113.740 14.855 ;
        RECT 113.930 14.685 114.100 14.855 ;
        RECT 114.290 14.685 114.460 14.855 ;
        RECT 114.650 14.685 114.820 14.855 ;
        RECT 115.010 14.685 115.180 14.855 ;
        RECT 115.370 14.685 115.540 14.855 ;
        RECT 115.730 14.685 115.900 14.855 ;
        RECT 116.090 14.685 116.260 14.855 ;
        RECT 116.450 14.685 116.620 14.855 ;
        RECT 116.810 14.685 116.980 14.855 ;
        RECT 117.170 14.685 117.340 14.855 ;
        RECT 117.530 14.685 117.700 14.855 ;
        RECT 117.890 14.685 118.060 14.855 ;
        RECT 56.330 13.540 56.500 13.710 ;
        RECT 56.690 13.540 56.860 13.710 ;
        RECT 57.050 13.540 57.220 13.710 ;
        RECT 57.410 13.540 57.580 13.710 ;
        RECT 57.770 13.540 57.940 13.710 ;
        RECT 58.130 13.540 58.300 13.710 ;
        RECT 58.490 13.540 58.660 13.710 ;
        RECT 58.850 13.540 59.020 13.710 ;
        RECT 59.210 13.540 59.380 13.710 ;
        RECT 59.570 13.540 59.740 13.710 ;
        RECT 59.930 13.540 60.100 13.710 ;
        RECT 60.290 13.540 60.460 13.710 ;
        RECT 60.650 13.540 60.820 13.710 ;
        RECT 61.010 13.540 61.180 13.710 ;
        RECT 61.370 13.540 61.540 13.710 ;
        RECT 61.730 13.540 61.900 13.710 ;
        RECT 62.090 13.540 62.260 13.710 ;
        RECT 62.450 13.540 62.620 13.710 ;
        RECT 62.810 13.540 62.980 13.710 ;
        RECT 63.170 13.540 63.340 13.710 ;
        RECT 63.530 13.540 63.700 13.710 ;
        RECT 63.890 13.540 64.060 13.710 ;
        RECT 64.250 13.540 64.420 13.710 ;
        RECT 64.610 13.540 64.780 13.710 ;
        RECT 64.970 13.540 65.140 13.710 ;
        RECT 65.330 13.540 65.500 13.710 ;
        RECT 65.690 13.540 65.860 13.710 ;
        RECT 66.050 13.540 66.220 13.710 ;
        RECT 66.410 13.540 66.580 13.710 ;
        RECT 66.770 13.540 66.940 13.710 ;
        RECT 67.130 13.540 67.300 13.710 ;
        RECT 67.490 13.540 67.660 13.710 ;
        RECT 67.850 13.540 68.020 13.710 ;
        RECT 68.210 13.540 68.380 13.710 ;
        RECT 68.570 13.540 68.740 13.710 ;
        RECT 68.930 13.540 69.100 13.710 ;
        RECT 69.290 13.540 69.460 13.710 ;
        RECT 69.650 13.540 69.820 13.710 ;
        RECT 70.010 13.540 70.180 13.710 ;
        RECT 70.370 13.540 70.540 13.710 ;
        RECT 70.730 13.540 70.900 13.710 ;
        RECT 71.090 13.540 71.260 13.710 ;
        RECT 71.450 13.540 71.620 13.710 ;
        RECT 71.810 13.540 71.980 13.710 ;
        RECT 72.170 13.540 72.340 13.710 ;
        RECT 72.530 13.540 72.700 13.710 ;
        RECT 72.890 13.540 73.060 13.710 ;
        RECT 73.250 13.540 73.420 13.710 ;
        RECT 73.610 13.540 73.780 13.710 ;
        RECT 73.970 13.540 74.140 13.710 ;
        RECT 74.330 13.540 74.500 13.710 ;
        RECT 74.690 13.540 74.860 13.710 ;
        RECT 75.050 13.540 75.220 13.710 ;
        RECT 75.410 13.540 75.580 13.710 ;
        RECT 75.770 13.540 75.940 13.710 ;
        RECT 76.130 13.540 76.300 13.710 ;
        RECT 76.490 13.540 76.660 13.710 ;
        RECT 76.850 13.540 77.020 13.710 ;
        RECT 77.210 13.540 77.380 13.710 ;
        RECT 77.570 13.540 77.740 13.710 ;
        RECT 77.930 13.540 78.100 13.710 ;
        RECT 78.290 13.540 78.460 13.710 ;
        RECT 78.650 13.540 78.820 13.710 ;
        RECT 79.010 13.540 79.180 13.710 ;
        RECT 79.370 13.540 79.540 13.710 ;
        RECT 79.730 13.540 79.900 13.710 ;
        RECT 80.090 13.540 80.260 13.710 ;
        RECT 80.450 13.540 80.620 13.710 ;
        RECT 80.810 13.540 80.980 13.710 ;
        RECT 81.170 13.540 81.340 13.710 ;
        RECT 81.530 13.540 81.700 13.710 ;
        RECT 81.890 13.540 82.060 13.710 ;
        RECT 82.250 13.540 82.420 13.710 ;
        RECT 82.610 13.540 82.780 13.710 ;
        RECT 82.970 13.540 83.140 13.710 ;
        RECT 83.330 13.540 83.500 13.710 ;
        RECT 83.690 13.540 83.860 13.710 ;
        RECT 84.050 13.540 84.220 13.710 ;
        RECT 84.410 13.540 84.580 13.710 ;
        RECT 84.770 13.540 84.940 13.710 ;
        RECT 85.130 13.540 85.300 13.710 ;
        RECT 85.490 13.540 85.660 13.710 ;
        RECT 85.850 13.540 86.020 13.710 ;
        RECT 86.210 13.540 86.380 13.710 ;
        RECT 86.570 13.540 86.740 13.710 ;
        RECT 86.930 13.540 87.100 13.710 ;
        RECT 87.290 13.540 87.460 13.710 ;
        RECT 87.650 13.540 87.820 13.710 ;
        RECT 88.010 13.540 88.180 13.710 ;
        RECT 88.370 13.540 88.540 13.710 ;
        RECT 88.730 13.540 88.900 13.710 ;
        RECT 89.090 13.540 89.260 13.710 ;
        RECT 89.450 13.540 89.620 13.710 ;
        RECT 89.810 13.540 89.980 13.710 ;
        RECT 90.170 13.540 90.340 13.710 ;
        RECT 90.530 13.540 90.700 13.710 ;
        RECT 90.890 13.540 91.060 13.710 ;
        RECT 91.250 13.540 91.420 13.710 ;
        RECT 91.610 13.540 91.780 13.710 ;
        RECT 91.970 13.540 92.140 13.710 ;
        RECT 92.330 13.540 92.500 13.710 ;
        RECT 92.690 13.540 92.860 13.710 ;
        RECT 93.050 13.540 93.220 13.710 ;
        RECT 93.410 13.540 93.580 13.710 ;
        RECT 93.770 13.540 93.940 13.710 ;
        RECT 94.130 13.540 94.300 13.710 ;
        RECT 94.490 13.540 94.660 13.710 ;
        RECT 94.850 13.540 95.020 13.710 ;
        RECT 55.980 13.240 56.150 13.410 ;
        RECT 95.480 13.240 95.650 13.410 ;
        RECT 55.980 12.880 56.150 13.050 ;
        RECT 58.630 12.990 58.800 13.160 ;
        RECT 58.990 12.990 59.160 13.160 ;
        RECT 59.350 12.990 59.520 13.160 ;
        RECT 59.710 12.990 59.880 13.160 ;
        RECT 60.070 12.990 60.240 13.160 ;
        RECT 60.910 12.990 61.080 13.160 ;
        RECT 61.270 12.990 61.440 13.160 ;
        RECT 61.630 12.990 61.800 13.160 ;
        RECT 61.990 12.990 62.160 13.160 ;
        RECT 62.350 12.990 62.520 13.160 ;
        RECT 66.310 12.990 66.480 13.160 ;
        RECT 66.670 12.990 66.840 13.160 ;
        RECT 67.030 12.990 67.200 13.160 ;
        RECT 67.390 12.990 67.560 13.160 ;
        RECT 67.750 12.990 67.920 13.160 ;
        RECT 68.590 12.990 68.760 13.160 ;
        RECT 68.950 12.990 69.120 13.160 ;
        RECT 69.310 12.990 69.480 13.160 ;
        RECT 69.670 12.990 69.840 13.160 ;
        RECT 70.030 12.990 70.200 13.160 ;
        RECT 70.870 12.990 71.040 13.160 ;
        RECT 71.230 12.990 71.400 13.160 ;
        RECT 71.590 12.990 71.760 13.160 ;
        RECT 71.950 12.990 72.120 13.160 ;
        RECT 72.310 12.990 72.480 13.160 ;
        RECT 73.150 12.990 73.320 13.160 ;
        RECT 73.510 12.990 73.680 13.160 ;
        RECT 73.870 12.990 74.040 13.160 ;
        RECT 74.230 12.990 74.400 13.160 ;
        RECT 74.590 12.990 74.760 13.160 ;
        RECT 75.430 12.990 75.600 13.160 ;
        RECT 75.790 12.990 75.960 13.160 ;
        RECT 76.150 12.990 76.320 13.160 ;
        RECT 76.510 12.990 76.680 13.160 ;
        RECT 76.870 12.990 77.040 13.160 ;
        RECT 77.710 12.990 77.880 13.160 ;
        RECT 78.070 12.990 78.240 13.160 ;
        RECT 78.430 12.990 78.600 13.160 ;
        RECT 78.790 12.990 78.960 13.160 ;
        RECT 79.150 12.990 79.320 13.160 ;
        RECT 79.990 12.990 80.160 13.160 ;
        RECT 80.350 12.990 80.520 13.160 ;
        RECT 80.710 12.990 80.880 13.160 ;
        RECT 81.070 12.990 81.240 13.160 ;
        RECT 81.430 12.990 81.600 13.160 ;
        RECT 82.270 12.990 82.440 13.160 ;
        RECT 82.630 12.990 82.800 13.160 ;
        RECT 82.990 12.990 83.160 13.160 ;
        RECT 83.350 12.990 83.520 13.160 ;
        RECT 83.710 12.990 83.880 13.160 ;
        RECT 84.550 12.990 84.720 13.160 ;
        RECT 84.910 12.990 85.080 13.160 ;
        RECT 85.270 12.990 85.440 13.160 ;
        RECT 85.630 12.990 85.800 13.160 ;
        RECT 85.990 12.990 86.160 13.160 ;
        RECT 86.830 12.990 87.000 13.160 ;
        RECT 87.190 12.990 87.360 13.160 ;
        RECT 87.550 12.990 87.720 13.160 ;
        RECT 87.910 12.990 88.080 13.160 ;
        RECT 88.270 12.990 88.440 13.160 ;
        RECT 89.110 12.990 89.280 13.160 ;
        RECT 89.470 12.990 89.640 13.160 ;
        RECT 89.830 12.990 90.000 13.160 ;
        RECT 90.190 12.990 90.360 13.160 ;
        RECT 90.550 12.990 90.720 13.160 ;
        RECT 91.390 12.990 91.560 13.160 ;
        RECT 91.750 12.990 91.920 13.160 ;
        RECT 92.110 12.990 92.280 13.160 ;
        RECT 92.470 12.990 92.640 13.160 ;
        RECT 92.830 12.990 93.000 13.160 ;
        RECT 95.480 12.880 95.650 13.050 ;
        RECT 55.980 12.520 56.150 12.690 ;
        RECT 55.980 12.160 56.150 12.330 ;
        RECT 55.980 11.800 56.150 11.970 ;
        RECT 56.650 12.335 56.820 12.505 ;
        RECT 56.650 11.975 56.820 12.145 ;
        RECT 57.430 12.335 57.600 12.505 ;
        RECT 57.430 11.975 57.600 12.145 ;
        RECT 58.210 12.335 58.380 12.505 ;
        RECT 58.210 11.975 58.380 12.145 ;
        RECT 60.490 12.335 60.660 12.505 ;
        RECT 60.490 11.975 60.660 12.145 ;
        RECT 62.770 12.335 62.940 12.505 ;
        RECT 62.770 11.975 62.940 12.145 ;
        RECT 63.550 12.335 63.720 12.505 ;
        RECT 63.550 11.975 63.720 12.145 ;
        RECT 64.330 12.335 64.500 12.505 ;
        RECT 64.330 11.975 64.500 12.145 ;
        RECT 65.110 12.335 65.280 12.505 ;
        RECT 65.110 11.975 65.280 12.145 ;
        RECT 65.890 12.335 66.060 12.505 ;
        RECT 65.890 11.975 66.060 12.145 ;
        RECT 68.170 12.335 68.340 12.505 ;
        RECT 68.170 11.975 68.340 12.145 ;
        RECT 70.450 12.335 70.620 12.505 ;
        RECT 70.450 11.975 70.620 12.145 ;
        RECT 72.730 12.335 72.900 12.505 ;
        RECT 72.730 11.975 72.900 12.145 ;
        RECT 75.010 12.335 75.180 12.505 ;
        RECT 75.010 11.975 75.180 12.145 ;
        RECT 77.290 12.335 77.460 12.505 ;
        RECT 77.290 11.975 77.460 12.145 ;
        RECT 79.570 12.335 79.740 12.505 ;
        RECT 79.570 11.975 79.740 12.145 ;
        RECT 81.850 12.335 82.020 12.505 ;
        RECT 81.850 11.975 82.020 12.145 ;
        RECT 84.130 12.335 84.300 12.505 ;
        RECT 84.130 11.975 84.300 12.145 ;
        RECT 86.410 12.335 86.580 12.505 ;
        RECT 86.410 11.975 86.580 12.145 ;
        RECT 88.690 12.335 88.860 12.505 ;
        RECT 88.690 11.975 88.860 12.145 ;
        RECT 90.970 12.335 91.140 12.505 ;
        RECT 90.970 11.975 91.140 12.145 ;
        RECT 93.250 12.335 93.420 12.505 ;
        RECT 93.250 11.975 93.420 12.145 ;
        RECT 94.030 12.335 94.200 12.505 ;
        RECT 94.030 11.975 94.200 12.145 ;
        RECT 94.810 12.335 94.980 12.505 ;
        RECT 94.810 11.975 94.980 12.145 ;
        RECT 95.480 12.520 95.650 12.690 ;
        RECT 95.480 12.160 95.650 12.330 ;
        RECT 95.480 11.800 95.650 11.970 ;
        RECT 55.980 11.440 56.150 11.610 ;
        RECT 55.980 11.080 56.150 11.250 ;
        RECT 57.070 11.320 57.240 11.490 ;
        RECT 57.430 11.320 57.600 11.490 ;
        RECT 57.790 11.320 57.960 11.490 ;
        RECT 63.190 11.320 63.360 11.490 ;
        RECT 63.550 11.320 63.720 11.490 ;
        RECT 63.910 11.320 64.080 11.490 ;
        RECT 64.750 11.320 64.920 11.490 ;
        RECT 65.110 11.320 65.280 11.490 ;
        RECT 65.470 11.320 65.640 11.490 ;
        RECT 66.310 11.320 66.480 11.490 ;
        RECT 66.670 11.320 66.840 11.490 ;
        RECT 67.030 11.320 67.200 11.490 ;
        RECT 67.390 11.320 67.560 11.490 ;
        RECT 67.750 11.320 67.920 11.490 ;
        RECT 68.590 11.320 68.760 11.490 ;
        RECT 68.950 11.320 69.120 11.490 ;
        RECT 69.310 11.320 69.480 11.490 ;
        RECT 69.670 11.320 69.840 11.490 ;
        RECT 70.030 11.320 70.200 11.490 ;
        RECT 70.870 11.320 71.040 11.490 ;
        RECT 71.230 11.320 71.400 11.490 ;
        RECT 71.590 11.320 71.760 11.490 ;
        RECT 71.950 11.320 72.120 11.490 ;
        RECT 72.310 11.320 72.480 11.490 ;
        RECT 73.150 11.320 73.320 11.490 ;
        RECT 73.510 11.320 73.680 11.490 ;
        RECT 73.870 11.320 74.040 11.490 ;
        RECT 74.230 11.320 74.400 11.490 ;
        RECT 74.590 11.320 74.760 11.490 ;
        RECT 75.430 11.320 75.600 11.490 ;
        RECT 75.790 11.320 75.960 11.490 ;
        RECT 76.150 11.320 76.320 11.490 ;
        RECT 76.510 11.320 76.680 11.490 ;
        RECT 76.870 11.320 77.040 11.490 ;
        RECT 77.710 11.320 77.880 11.490 ;
        RECT 78.070 11.320 78.240 11.490 ;
        RECT 78.430 11.320 78.600 11.490 ;
        RECT 78.790 11.320 78.960 11.490 ;
        RECT 79.150 11.320 79.320 11.490 ;
        RECT 79.990 11.320 80.160 11.490 ;
        RECT 80.350 11.320 80.520 11.490 ;
        RECT 80.710 11.320 80.880 11.490 ;
        RECT 81.070 11.320 81.240 11.490 ;
        RECT 81.430 11.320 81.600 11.490 ;
        RECT 82.270 11.320 82.440 11.490 ;
        RECT 82.630 11.320 82.800 11.490 ;
        RECT 82.990 11.320 83.160 11.490 ;
        RECT 83.350 11.320 83.520 11.490 ;
        RECT 83.710 11.320 83.880 11.490 ;
        RECT 84.550 11.320 84.720 11.490 ;
        RECT 84.910 11.320 85.080 11.490 ;
        RECT 85.270 11.320 85.440 11.490 ;
        RECT 85.630 11.320 85.800 11.490 ;
        RECT 85.990 11.320 86.160 11.490 ;
        RECT 86.830 11.320 87.000 11.490 ;
        RECT 87.190 11.320 87.360 11.490 ;
        RECT 87.550 11.320 87.720 11.490 ;
        RECT 87.910 11.320 88.080 11.490 ;
        RECT 88.270 11.320 88.440 11.490 ;
        RECT 89.110 11.320 89.280 11.490 ;
        RECT 89.470 11.320 89.640 11.490 ;
        RECT 89.830 11.320 90.000 11.490 ;
        RECT 90.190 11.320 90.360 11.490 ;
        RECT 90.550 11.320 90.720 11.490 ;
        RECT 91.390 11.320 91.560 11.490 ;
        RECT 91.750 11.320 91.920 11.490 ;
        RECT 92.110 11.320 92.280 11.490 ;
        RECT 92.470 11.320 92.640 11.490 ;
        RECT 92.830 11.320 93.000 11.490 ;
        RECT 93.670 11.320 93.840 11.490 ;
        RECT 94.030 11.320 94.200 11.490 ;
        RECT 94.390 11.320 94.560 11.490 ;
        RECT 95.480 11.440 95.650 11.610 ;
        RECT 55.980 10.720 56.150 10.890 ;
        RECT 55.980 10.360 56.150 10.530 ;
        RECT 55.980 10.000 56.150 10.170 ;
        RECT 55.980 9.640 56.150 9.810 ;
        RECT 95.480 11.080 95.650 11.250 ;
        RECT 95.480 10.720 95.650 10.890 ;
        RECT 95.480 10.360 95.650 10.530 ;
        RECT 95.480 10.000 95.650 10.170 ;
        RECT 55.980 9.280 56.150 9.450 ;
        RECT 66.310 9.400 66.480 9.570 ;
        RECT 66.670 9.400 66.840 9.570 ;
        RECT 67.030 9.400 67.200 9.570 ;
        RECT 67.390 9.400 67.560 9.570 ;
        RECT 67.750 9.400 67.920 9.570 ;
        RECT 68.590 9.400 68.760 9.570 ;
        RECT 68.950 9.400 69.120 9.570 ;
        RECT 69.310 9.400 69.480 9.570 ;
        RECT 69.670 9.400 69.840 9.570 ;
        RECT 70.030 9.400 70.200 9.570 ;
        RECT 70.870 9.400 71.040 9.570 ;
        RECT 71.230 9.400 71.400 9.570 ;
        RECT 71.590 9.400 71.760 9.570 ;
        RECT 71.950 9.400 72.120 9.570 ;
        RECT 72.310 9.400 72.480 9.570 ;
        RECT 73.150 9.400 73.320 9.570 ;
        RECT 73.510 9.400 73.680 9.570 ;
        RECT 73.870 9.400 74.040 9.570 ;
        RECT 74.230 9.400 74.400 9.570 ;
        RECT 74.590 9.400 74.760 9.570 ;
        RECT 75.430 9.400 75.600 9.570 ;
        RECT 75.790 9.400 75.960 9.570 ;
        RECT 76.150 9.400 76.320 9.570 ;
        RECT 76.510 9.400 76.680 9.570 ;
        RECT 76.870 9.400 77.040 9.570 ;
        RECT 82.270 9.400 82.440 9.570 ;
        RECT 82.630 9.400 82.800 9.570 ;
        RECT 82.990 9.400 83.160 9.570 ;
        RECT 83.350 9.400 83.520 9.570 ;
        RECT 83.710 9.400 83.880 9.570 ;
        RECT 84.550 9.400 84.720 9.570 ;
        RECT 84.910 9.400 85.080 9.570 ;
        RECT 85.270 9.400 85.440 9.570 ;
        RECT 85.630 9.400 85.800 9.570 ;
        RECT 85.990 9.400 86.160 9.570 ;
        RECT 86.830 9.400 87.000 9.570 ;
        RECT 87.190 9.400 87.360 9.570 ;
        RECT 87.550 9.400 87.720 9.570 ;
        RECT 87.910 9.400 88.080 9.570 ;
        RECT 88.270 9.400 88.440 9.570 ;
        RECT 89.110 9.400 89.280 9.570 ;
        RECT 89.470 9.400 89.640 9.570 ;
        RECT 89.830 9.400 90.000 9.570 ;
        RECT 90.190 9.400 90.360 9.570 ;
        RECT 90.550 9.400 90.720 9.570 ;
        RECT 91.390 9.400 91.560 9.570 ;
        RECT 91.750 9.400 91.920 9.570 ;
        RECT 92.110 9.400 92.280 9.570 ;
        RECT 92.470 9.400 92.640 9.570 ;
        RECT 92.830 9.400 93.000 9.570 ;
        RECT 95.480 9.640 95.650 9.810 ;
        RECT 95.480 9.280 95.650 9.450 ;
        RECT 55.980 8.920 56.150 9.090 ;
        RECT 55.980 8.560 56.150 8.730 ;
        RECT 55.980 8.200 56.150 8.370 ;
        RECT 65.890 8.745 66.060 8.915 ;
        RECT 65.890 8.385 66.060 8.555 ;
        RECT 68.170 8.745 68.340 8.915 ;
        RECT 68.170 8.385 68.340 8.555 ;
        RECT 70.450 8.745 70.620 8.915 ;
        RECT 70.450 8.385 70.620 8.555 ;
        RECT 72.730 8.745 72.900 8.915 ;
        RECT 72.730 8.385 72.900 8.555 ;
        RECT 75.010 8.745 75.180 8.915 ;
        RECT 75.010 8.385 75.180 8.555 ;
        RECT 77.290 8.745 77.460 8.915 ;
        RECT 77.290 8.385 77.460 8.555 ;
        RECT 79.570 8.745 79.740 8.915 ;
        RECT 79.570 8.385 79.740 8.555 ;
        RECT 81.850 8.745 82.020 8.915 ;
        RECT 81.850 8.385 82.020 8.555 ;
        RECT 84.130 8.745 84.300 8.915 ;
        RECT 84.130 8.385 84.300 8.555 ;
        RECT 86.410 8.745 86.580 8.915 ;
        RECT 86.410 8.385 86.580 8.555 ;
        RECT 88.690 8.745 88.860 8.915 ;
        RECT 88.690 8.385 88.860 8.555 ;
        RECT 90.970 8.745 91.140 8.915 ;
        RECT 90.970 8.385 91.140 8.555 ;
        RECT 93.250 8.745 93.420 8.915 ;
        RECT 93.250 8.385 93.420 8.555 ;
        RECT 95.480 8.920 95.650 9.090 ;
        RECT 95.480 8.560 95.650 8.730 ;
        RECT 95.480 8.200 95.650 8.370 ;
        RECT 55.980 7.840 56.150 8.010 ;
        RECT 77.710 7.730 77.880 7.900 ;
        RECT 78.070 7.730 78.240 7.900 ;
        RECT 78.430 7.730 78.600 7.900 ;
        RECT 78.790 7.730 78.960 7.900 ;
        RECT 79.150 7.730 79.320 7.900 ;
        RECT 79.990 7.730 80.160 7.900 ;
        RECT 80.350 7.730 80.520 7.900 ;
        RECT 80.710 7.730 80.880 7.900 ;
        RECT 81.070 7.730 81.240 7.900 ;
        RECT 81.430 7.730 81.600 7.900 ;
        RECT 95.480 7.840 95.650 8.010 ;
        RECT 55.980 7.480 56.150 7.650 ;
        RECT 95.480 7.480 95.650 7.650 ;
        RECT 56.330 7.180 56.500 7.350 ;
        RECT 56.690 7.180 56.860 7.350 ;
        RECT 57.050 7.180 57.220 7.350 ;
        RECT 57.410 7.180 57.580 7.350 ;
        RECT 57.770 7.180 57.940 7.350 ;
        RECT 58.130 7.180 58.300 7.350 ;
        RECT 58.490 7.180 58.660 7.350 ;
        RECT 58.850 7.180 59.020 7.350 ;
        RECT 59.210 7.180 59.380 7.350 ;
        RECT 59.570 7.180 59.740 7.350 ;
        RECT 59.930 7.180 60.100 7.350 ;
        RECT 60.290 7.180 60.460 7.350 ;
        RECT 60.650 7.180 60.820 7.350 ;
        RECT 61.010 7.180 61.180 7.350 ;
        RECT 61.370 7.180 61.540 7.350 ;
        RECT 61.730 7.180 61.900 7.350 ;
        RECT 62.090 7.180 62.260 7.350 ;
        RECT 62.450 7.180 62.620 7.350 ;
        RECT 62.810 7.180 62.980 7.350 ;
        RECT 63.170 7.180 63.340 7.350 ;
        RECT 63.530 7.180 63.700 7.350 ;
        RECT 63.890 7.180 64.060 7.350 ;
        RECT 64.250 7.180 64.420 7.350 ;
        RECT 64.610 7.180 64.780 7.350 ;
        RECT 64.970 7.180 65.140 7.350 ;
        RECT 65.330 7.180 65.500 7.350 ;
        RECT 65.690 7.180 65.860 7.350 ;
        RECT 66.050 7.180 66.220 7.350 ;
        RECT 66.410 7.180 66.580 7.350 ;
        RECT 66.770 7.180 66.940 7.350 ;
        RECT 67.130 7.180 67.300 7.350 ;
        RECT 67.490 7.180 67.660 7.350 ;
        RECT 67.850 7.180 68.020 7.350 ;
        RECT 68.210 7.180 68.380 7.350 ;
        RECT 68.570 7.180 68.740 7.350 ;
        RECT 68.930 7.180 69.100 7.350 ;
        RECT 69.290 7.180 69.460 7.350 ;
        RECT 69.650 7.180 69.820 7.350 ;
        RECT 70.010 7.180 70.180 7.350 ;
        RECT 70.370 7.180 70.540 7.350 ;
        RECT 70.730 7.180 70.900 7.350 ;
        RECT 71.090 7.180 71.260 7.350 ;
        RECT 71.450 7.180 71.620 7.350 ;
        RECT 71.810 7.180 71.980 7.350 ;
        RECT 72.170 7.180 72.340 7.350 ;
        RECT 72.530 7.180 72.700 7.350 ;
        RECT 72.890 7.180 73.060 7.350 ;
        RECT 73.250 7.180 73.420 7.350 ;
        RECT 73.610 7.180 73.780 7.350 ;
        RECT 73.970 7.180 74.140 7.350 ;
        RECT 74.330 7.180 74.500 7.350 ;
        RECT 74.690 7.180 74.860 7.350 ;
        RECT 75.050 7.180 75.220 7.350 ;
        RECT 75.410 7.180 75.580 7.350 ;
        RECT 75.770 7.180 75.940 7.350 ;
        RECT 76.130 7.180 76.300 7.350 ;
        RECT 76.490 7.180 76.660 7.350 ;
        RECT 76.850 7.180 77.020 7.350 ;
        RECT 77.210 7.180 77.380 7.350 ;
        RECT 77.570 7.180 77.740 7.350 ;
        RECT 77.930 7.180 78.100 7.350 ;
        RECT 78.290 7.180 78.460 7.350 ;
        RECT 78.650 7.180 78.820 7.350 ;
        RECT 79.010 7.180 79.180 7.350 ;
        RECT 79.370 7.180 79.540 7.350 ;
        RECT 79.730 7.180 79.900 7.350 ;
        RECT 80.090 7.180 80.260 7.350 ;
        RECT 80.450 7.180 80.620 7.350 ;
        RECT 80.810 7.180 80.980 7.350 ;
        RECT 81.170 7.180 81.340 7.350 ;
        RECT 81.530 7.180 81.700 7.350 ;
        RECT 81.890 7.180 82.060 7.350 ;
        RECT 82.250 7.180 82.420 7.350 ;
        RECT 82.610 7.180 82.780 7.350 ;
        RECT 82.970 7.180 83.140 7.350 ;
        RECT 83.330 7.180 83.500 7.350 ;
        RECT 83.690 7.180 83.860 7.350 ;
        RECT 84.050 7.180 84.220 7.350 ;
        RECT 84.410 7.180 84.580 7.350 ;
        RECT 84.770 7.180 84.940 7.350 ;
        RECT 85.130 7.180 85.300 7.350 ;
        RECT 85.490 7.180 85.660 7.350 ;
        RECT 85.850 7.180 86.020 7.350 ;
        RECT 86.210 7.180 86.380 7.350 ;
        RECT 86.570 7.180 86.740 7.350 ;
        RECT 86.930 7.180 87.100 7.350 ;
        RECT 87.290 7.180 87.460 7.350 ;
        RECT 87.650 7.180 87.820 7.350 ;
        RECT 88.010 7.180 88.180 7.350 ;
        RECT 88.370 7.180 88.540 7.350 ;
        RECT 88.730 7.180 88.900 7.350 ;
        RECT 89.090 7.180 89.260 7.350 ;
        RECT 89.450 7.180 89.620 7.350 ;
        RECT 89.810 7.180 89.980 7.350 ;
        RECT 90.170 7.180 90.340 7.350 ;
        RECT 90.530 7.180 90.700 7.350 ;
        RECT 90.890 7.180 91.060 7.350 ;
        RECT 91.250 7.180 91.420 7.350 ;
        RECT 91.610 7.180 91.780 7.350 ;
        RECT 91.970 7.180 92.140 7.350 ;
        RECT 92.330 7.180 92.500 7.350 ;
        RECT 92.690 7.180 92.860 7.350 ;
        RECT 93.050 7.180 93.220 7.350 ;
        RECT 93.410 7.180 93.580 7.350 ;
        RECT 93.770 7.180 93.940 7.350 ;
        RECT 94.130 7.180 94.300 7.350 ;
        RECT 94.490 7.180 94.660 7.350 ;
        RECT 94.850 7.180 95.020 7.350 ;
      LAYER met1 ;
        RECT 137.110 77.865 147.260 78.155 ;
        RECT 42.710 76.620 130.900 76.910 ;
        RECT 42.710 76.360 43.000 76.620 ;
        RECT 130.610 76.360 130.900 76.620 ;
        RECT 42.710 76.070 47.740 76.360 ;
        RECT 48.350 76.070 50.020 76.360 ;
        RECT 50.630 76.070 52.300 76.360 ;
        RECT 52.910 76.070 54.580 76.360 ;
        RECT 55.190 76.070 56.860 76.360 ;
        RECT 57.470 76.070 59.140 76.360 ;
        RECT 59.750 76.070 61.420 76.360 ;
        RECT 62.030 76.070 63.700 76.360 ;
        RECT 64.310 76.070 65.980 76.360 ;
        RECT 66.590 76.070 68.260 76.360 ;
        RECT 68.870 76.070 70.540 76.360 ;
        RECT 71.150 76.070 72.820 76.360 ;
        RECT 73.430 76.070 75.100 76.360 ;
        RECT 75.710 76.070 77.380 76.360 ;
        RECT 77.990 76.070 79.660 76.360 ;
        RECT 80.270 76.070 81.940 76.360 ;
        RECT 82.550 76.070 84.220 76.360 ;
        RECT 84.830 76.070 86.500 76.360 ;
        RECT 87.110 76.070 88.780 76.360 ;
        RECT 89.390 76.070 91.060 76.360 ;
        RECT 91.670 76.070 93.340 76.360 ;
        RECT 93.950 76.070 95.620 76.360 ;
        RECT 96.230 76.070 97.900 76.360 ;
        RECT 98.510 76.070 100.180 76.360 ;
        RECT 100.790 76.070 102.460 76.360 ;
        RECT 103.070 76.070 104.740 76.360 ;
        RECT 105.350 76.070 107.020 76.360 ;
        RECT 107.630 76.070 109.300 76.360 ;
        RECT 109.910 76.070 111.580 76.360 ;
        RECT 112.190 76.070 113.860 76.360 ;
        RECT 114.470 76.070 116.140 76.360 ;
        RECT 116.750 76.070 130.900 76.360 ;
        RECT 42.710 73.620 43.000 76.070 ;
        RECT 118.610 75.880 118.840 76.070 ;
        RECT 120.890 75.880 121.120 76.070 ;
        RECT 123.170 75.880 123.400 76.070 ;
        RECT 125.450 75.880 125.680 76.070 ;
        RECT 43.355 75.180 43.615 75.880 ;
        RECT 45.635 75.180 45.895 75.880 ;
        RECT 47.915 75.180 48.175 75.880 ;
        RECT 50.195 75.180 50.455 75.880 ;
        RECT 52.475 75.180 52.735 75.880 ;
        RECT 54.755 75.180 55.015 75.880 ;
        RECT 57.035 75.180 57.295 75.880 ;
        RECT 59.315 75.180 59.575 75.880 ;
        RECT 61.595 75.180 61.855 75.880 ;
        RECT 63.875 75.180 64.135 75.880 ;
        RECT 66.155 75.180 66.415 75.880 ;
        RECT 68.435 75.180 68.695 75.880 ;
        RECT 70.715 75.180 70.975 75.880 ;
        RECT 72.995 75.180 73.255 75.880 ;
        RECT 75.275 75.180 75.535 75.880 ;
        RECT 77.555 75.180 77.815 75.880 ;
        RECT 79.835 75.180 80.095 75.880 ;
        RECT 82.115 75.180 82.375 75.880 ;
        RECT 84.395 75.180 84.655 75.880 ;
        RECT 86.675 75.180 86.935 75.880 ;
        RECT 88.955 75.180 89.215 75.880 ;
        RECT 91.235 75.180 91.495 75.880 ;
        RECT 93.515 75.180 93.775 75.880 ;
        RECT 95.795 75.180 96.055 75.880 ;
        RECT 98.075 75.180 98.335 75.880 ;
        RECT 100.355 75.180 100.615 75.880 ;
        RECT 102.635 75.180 102.895 75.880 ;
        RECT 104.915 75.180 105.175 75.880 ;
        RECT 107.195 75.180 107.455 75.880 ;
        RECT 109.475 75.180 109.735 75.880 ;
        RECT 111.755 75.180 112.015 75.880 ;
        RECT 114.035 75.180 114.295 75.880 ;
        RECT 116.315 75.180 116.575 75.880 ;
        RECT 118.595 75.180 118.855 75.880 ;
        RECT 120.875 75.180 121.135 75.880 ;
        RECT 123.155 75.180 123.415 75.880 ;
        RECT 125.435 75.180 125.695 75.880 ;
        RECT 127.715 75.180 127.975 75.880 ;
        RECT 129.995 75.180 130.255 75.880 ;
        RECT 43.490 74.680 124.880 75.010 ;
        RECT 130.610 74.990 130.900 76.070 ;
        RECT 137.110 76.235 137.400 77.865 ;
        RECT 141.640 77.315 142.730 77.610 ;
        RECT 137.755 76.425 138.015 77.125 ;
        RECT 138.185 76.425 138.445 77.125 ;
        RECT 138.615 76.425 138.875 77.125 ;
        RECT 139.045 76.425 139.305 77.125 ;
        RECT 139.475 76.425 139.735 77.125 ;
        RECT 139.905 76.425 140.165 77.125 ;
        RECT 140.335 76.425 140.595 77.125 ;
        RECT 140.765 76.425 141.025 77.125 ;
        RECT 141.195 76.425 141.455 77.125 ;
        RECT 141.625 76.425 141.885 77.125 ;
        RECT 142.055 76.425 142.315 77.125 ;
        RECT 142.485 76.425 142.745 77.125 ;
        RECT 142.915 76.425 143.175 77.125 ;
        RECT 143.345 76.425 143.605 77.125 ;
        RECT 143.775 76.425 144.035 77.125 ;
        RECT 144.205 76.425 144.465 77.125 ;
        RECT 144.635 76.425 144.895 77.125 ;
        RECT 145.065 76.425 145.325 77.125 ;
        RECT 145.495 76.425 145.755 77.125 ;
        RECT 145.925 76.425 146.185 77.125 ;
        RECT 146.355 76.425 146.615 77.125 ;
        RECT 146.970 76.235 147.260 77.865 ;
        RECT 137.110 75.945 141.010 76.235 ;
        RECT 143.360 75.945 147.260 76.235 ;
        RECT 137.110 75.685 137.400 75.945 ;
        RECT 146.970 75.685 147.260 75.945 ;
        RECT 137.110 75.395 147.260 75.685 ;
        RECT 128.150 74.700 130.900 74.990 ;
        RECT 144.285 74.885 145.425 75.395 ;
        RECT 43.355 73.810 43.615 74.510 ;
        RECT 45.635 73.810 45.895 74.510 ;
        RECT 47.915 73.810 48.175 74.510 ;
        RECT 50.195 73.810 50.455 74.510 ;
        RECT 52.475 73.810 52.735 74.510 ;
        RECT 54.755 73.810 55.015 74.510 ;
        RECT 57.035 73.810 57.295 74.510 ;
        RECT 59.315 73.810 59.575 74.510 ;
        RECT 61.595 73.810 61.855 74.510 ;
        RECT 63.875 73.810 64.135 74.510 ;
        RECT 66.155 73.810 66.415 74.510 ;
        RECT 68.435 73.810 68.695 74.510 ;
        RECT 70.715 73.810 70.975 74.510 ;
        RECT 72.995 73.810 73.255 74.510 ;
        RECT 75.275 73.810 75.535 74.510 ;
        RECT 77.555 73.810 77.815 74.510 ;
        RECT 79.835 73.810 80.095 74.510 ;
        RECT 82.115 73.810 82.375 74.510 ;
        RECT 84.395 73.810 84.655 74.510 ;
        RECT 86.675 73.810 86.935 74.510 ;
        RECT 88.955 73.810 89.215 74.510 ;
        RECT 91.235 73.810 91.495 74.510 ;
        RECT 93.515 73.810 93.775 74.510 ;
        RECT 95.795 73.810 96.055 74.510 ;
        RECT 98.075 73.810 98.335 74.510 ;
        RECT 100.355 73.810 100.615 74.510 ;
        RECT 102.635 73.810 102.895 74.510 ;
        RECT 104.915 73.810 105.175 74.510 ;
        RECT 107.195 73.810 107.455 74.510 ;
        RECT 109.475 73.810 109.735 74.510 ;
        RECT 111.755 73.810 112.015 74.510 ;
        RECT 114.035 73.810 114.295 74.510 ;
        RECT 116.315 73.810 116.575 74.510 ;
        RECT 118.595 73.810 118.855 74.510 ;
        RECT 120.875 73.810 121.135 74.510 ;
        RECT 123.155 73.810 123.415 74.510 ;
        RECT 125.435 73.810 125.695 74.510 ;
        RECT 127.715 73.810 127.975 74.510 ;
        RECT 129.995 73.810 130.255 74.510 ;
        RECT 118.610 73.620 118.840 73.810 ;
        RECT 120.890 73.620 121.120 73.810 ;
        RECT 130.610 73.620 130.900 74.700 ;
        RECT 42.710 73.330 47.740 73.620 ;
        RECT 48.350 73.330 50.020 73.620 ;
        RECT 50.630 73.330 52.300 73.620 ;
        RECT 52.910 73.330 54.580 73.620 ;
        RECT 55.190 73.330 56.860 73.620 ;
        RECT 57.470 73.330 59.140 73.620 ;
        RECT 59.750 73.330 61.420 73.620 ;
        RECT 62.030 73.330 63.700 73.620 ;
        RECT 64.310 73.330 65.980 73.620 ;
        RECT 66.590 73.330 68.260 73.620 ;
        RECT 68.870 73.330 70.540 73.620 ;
        RECT 71.150 73.330 72.820 73.620 ;
        RECT 73.430 73.330 75.100 73.620 ;
        RECT 75.710 73.330 77.380 73.620 ;
        RECT 77.990 73.330 79.660 73.620 ;
        RECT 80.270 73.330 81.940 73.620 ;
        RECT 82.550 73.330 84.220 73.620 ;
        RECT 84.830 73.330 86.500 73.620 ;
        RECT 87.110 73.330 88.780 73.620 ;
        RECT 89.390 73.330 91.060 73.620 ;
        RECT 91.670 73.330 93.340 73.620 ;
        RECT 93.950 73.330 95.620 73.620 ;
        RECT 96.230 73.330 97.900 73.620 ;
        RECT 98.510 73.330 100.180 73.620 ;
        RECT 100.790 73.330 102.460 73.620 ;
        RECT 103.070 73.330 104.740 73.620 ;
        RECT 105.350 73.330 107.020 73.620 ;
        RECT 107.630 73.330 109.300 73.620 ;
        RECT 109.910 73.330 111.580 73.620 ;
        RECT 112.190 73.330 113.860 73.620 ;
        RECT 114.470 73.330 116.140 73.620 ;
        RECT 116.750 73.330 122.980 73.620 ;
        RECT 123.590 73.330 127.540 73.620 ;
        RECT 128.150 73.330 130.900 73.620 ;
        RECT 42.710 73.070 43.000 73.330 ;
        RECT 130.610 73.070 130.900 73.330 ;
        RECT 42.710 72.780 130.900 73.070 ;
        RECT 137.070 74.595 142.140 74.885 ;
        RECT 137.070 73.650 137.360 74.595 ;
        RECT 137.595 74.045 140.150 74.375 ;
        RECT 137.770 73.650 138.000 73.855 ;
        RECT 138.200 73.650 138.430 73.855 ;
        RECT 137.070 73.360 138.430 73.650 ;
        RECT 137.070 72.965 137.360 73.360 ;
        RECT 137.770 73.155 138.000 73.360 ;
        RECT 138.200 73.155 138.430 73.360 ;
        RECT 138.615 73.155 138.875 73.855 ;
        RECT 139.045 73.155 139.305 73.855 ;
        RECT 139.475 73.155 139.735 73.855 ;
        RECT 139.905 73.155 140.165 73.855 ;
        RECT 140.335 73.155 140.595 73.855 ;
        RECT 140.780 73.650 141.010 73.855 ;
        RECT 141.210 73.650 141.440 73.855 ;
        RECT 141.850 73.650 142.140 74.595 ;
        RECT 140.780 73.360 142.140 73.650 ;
        RECT 140.780 73.155 141.010 73.360 ;
        RECT 141.210 73.155 141.440 73.360 ;
        RECT 141.850 72.965 142.140 73.360 ;
        RECT 92.215 72.195 94.215 72.780 ;
        RECT 128.215 72.195 130.215 72.780 ;
        RECT 137.070 72.675 138.430 72.965 ;
        RECT 140.780 72.675 142.140 72.965 ;
        RECT 89.500 71.905 97.930 72.195 ;
        RECT 89.500 70.775 89.790 71.905 ;
        RECT 93.165 71.355 94.260 71.685 ;
        RECT 90.160 70.775 90.390 71.165 ;
        RECT 90.590 70.775 90.820 71.165 ;
        RECT 91.020 70.775 91.250 71.165 ;
        RECT 91.450 70.775 91.680 71.165 ;
        RECT 91.880 70.775 92.110 71.165 ;
        RECT 92.310 70.775 92.540 71.165 ;
        RECT 92.740 70.775 92.970 71.165 ;
        RECT 89.500 70.485 92.970 70.775 ;
        RECT 89.500 69.975 89.790 70.485 ;
        RECT 90.160 70.165 90.390 70.485 ;
        RECT 90.590 70.165 90.820 70.485 ;
        RECT 91.020 70.165 91.250 70.485 ;
        RECT 91.450 70.165 91.680 70.485 ;
        RECT 91.880 70.165 92.110 70.485 ;
        RECT 92.310 70.165 92.540 70.485 ;
        RECT 92.740 70.165 92.970 70.485 ;
        RECT 93.155 70.165 93.415 71.165 ;
        RECT 89.500 69.685 92.540 69.975 ;
        RECT 89.500 69.425 89.790 69.685 ;
        RECT 93.600 69.425 93.830 71.165 ;
        RECT 94.015 70.165 94.275 71.165 ;
        RECT 94.460 70.775 94.690 71.165 ;
        RECT 94.890 70.775 95.120 71.165 ;
        RECT 95.320 70.775 95.550 71.165 ;
        RECT 95.750 70.775 95.980 71.165 ;
        RECT 96.180 70.775 96.410 71.165 ;
        RECT 96.610 70.775 96.840 71.165 ;
        RECT 97.040 70.775 97.270 71.165 ;
        RECT 97.640 70.775 97.930 71.905 ;
        RECT 94.460 70.485 97.930 70.775 ;
        RECT 94.460 70.165 94.690 70.485 ;
        RECT 94.890 70.165 95.120 70.485 ;
        RECT 95.320 70.165 95.550 70.485 ;
        RECT 95.750 70.165 95.980 70.485 ;
        RECT 96.180 70.165 96.410 70.485 ;
        RECT 96.610 70.165 96.840 70.485 ;
        RECT 97.040 70.165 97.270 70.485 ;
        RECT 97.640 69.975 97.930 70.485 ;
        RECT 94.890 69.685 97.930 69.975 ;
        RECT 97.640 69.425 97.930 69.685 ;
        RECT 89.500 69.135 97.930 69.425 ;
        RECT 123.700 71.905 132.130 72.195 ;
        RECT 123.700 70.775 123.990 71.905 ;
        RECT 127.365 71.355 128.460 71.685 ;
        RECT 124.360 70.775 124.590 71.165 ;
        RECT 124.790 70.775 125.020 71.165 ;
        RECT 125.220 70.775 125.450 71.165 ;
        RECT 125.650 70.775 125.880 71.165 ;
        RECT 126.080 70.775 126.310 71.165 ;
        RECT 126.510 70.775 126.740 71.165 ;
        RECT 126.940 70.775 127.170 71.165 ;
        RECT 123.700 70.485 127.170 70.775 ;
        RECT 123.700 69.975 123.990 70.485 ;
        RECT 124.360 70.165 124.590 70.485 ;
        RECT 124.790 70.165 125.020 70.485 ;
        RECT 125.220 70.165 125.450 70.485 ;
        RECT 125.650 70.165 125.880 70.485 ;
        RECT 126.080 70.165 126.310 70.485 ;
        RECT 126.510 70.165 126.740 70.485 ;
        RECT 126.940 70.165 127.170 70.485 ;
        RECT 127.355 70.165 127.615 71.165 ;
        RECT 123.700 69.685 126.740 69.975 ;
        RECT 123.700 69.425 123.990 69.685 ;
        RECT 127.800 69.425 128.030 71.165 ;
        RECT 128.215 70.165 128.475 71.165 ;
        RECT 128.660 70.775 128.890 71.165 ;
        RECT 129.090 70.775 129.320 71.165 ;
        RECT 129.520 70.775 129.750 71.165 ;
        RECT 129.950 70.775 130.180 71.165 ;
        RECT 130.380 70.775 130.610 71.165 ;
        RECT 130.810 70.775 131.040 71.165 ;
        RECT 131.240 70.775 131.470 71.165 ;
        RECT 131.840 70.775 132.130 71.905 ;
        RECT 128.660 70.485 132.130 70.775 ;
        RECT 128.660 70.165 128.890 70.485 ;
        RECT 129.090 70.165 129.320 70.485 ;
        RECT 129.520 70.165 129.750 70.485 ;
        RECT 129.950 70.165 130.180 70.485 ;
        RECT 130.380 70.165 130.610 70.485 ;
        RECT 130.810 70.165 131.040 70.485 ;
        RECT 131.240 70.165 131.470 70.485 ;
        RECT 131.840 69.975 132.130 70.485 ;
        RECT 129.090 69.685 132.130 69.975 ;
        RECT 131.840 69.425 132.130 69.685 ;
        RECT 123.700 69.135 132.130 69.425 ;
        RECT 137.070 70.250 137.360 72.675 ;
        RECT 137.670 71.330 140.150 71.660 ;
        RECT 137.755 70.440 138.015 71.140 ;
        RECT 138.185 70.440 138.445 71.140 ;
        RECT 138.615 70.440 138.875 71.140 ;
        RECT 139.030 70.440 139.290 71.140 ;
        RECT 139.475 70.440 139.735 71.140 ;
        RECT 139.890 70.440 140.150 71.140 ;
        RECT 140.335 70.440 140.595 71.140 ;
        RECT 140.765 70.440 141.025 71.140 ;
        RECT 141.195 70.440 141.455 71.140 ;
        RECT 141.850 70.250 142.140 72.675 ;
        RECT 137.070 69.960 138.430 70.250 ;
        RECT 140.780 69.960 142.140 70.250 ;
        RECT 137.070 69.700 137.360 69.960 ;
        RECT 141.850 69.700 142.140 69.960 ;
        RECT 137.070 69.410 142.140 69.700 ;
        RECT 142.360 74.595 147.350 74.885 ;
        RECT 142.360 73.650 142.650 74.595 ;
        RECT 144.310 74.045 146.715 74.375 ;
        RECT 143.020 73.650 143.250 73.855 ;
        RECT 143.450 73.650 143.680 73.855 ;
        RECT 142.360 73.360 143.680 73.650 ;
        RECT 142.360 72.965 142.650 73.360 ;
        RECT 143.020 73.155 143.250 73.360 ;
        RECT 143.450 73.155 143.680 73.360 ;
        RECT 143.865 73.155 144.125 73.855 ;
        RECT 144.295 73.155 144.555 73.855 ;
        RECT 144.725 73.155 144.985 73.855 ;
        RECT 145.155 73.155 145.415 73.855 ;
        RECT 145.585 73.155 145.845 73.855 ;
        RECT 146.030 73.650 146.260 73.855 ;
        RECT 146.460 73.650 146.690 73.855 ;
        RECT 147.060 73.650 147.350 74.595 ;
        RECT 146.030 73.360 147.350 73.650 ;
        RECT 146.030 73.155 146.260 73.360 ;
        RECT 146.460 73.155 146.690 73.360 ;
        RECT 147.060 72.965 147.350 73.360 ;
        RECT 142.360 72.675 143.680 72.965 ;
        RECT 146.030 72.675 147.350 72.965 ;
        RECT 142.360 70.250 142.650 72.675 ;
        RECT 142.935 71.660 144.025 71.770 ;
        RECT 142.935 71.330 145.400 71.660 ;
        RECT 143.005 70.440 143.265 71.140 ;
        RECT 143.435 70.440 143.695 71.140 ;
        RECT 143.865 70.440 144.125 71.140 ;
        RECT 144.280 70.440 144.540 71.140 ;
        RECT 144.725 70.440 144.985 71.140 ;
        RECT 145.140 70.440 145.400 71.140 ;
        RECT 145.585 70.440 145.845 71.140 ;
        RECT 146.015 70.440 146.275 71.140 ;
        RECT 146.445 70.440 146.705 71.140 ;
        RECT 147.060 70.250 147.350 72.675 ;
        RECT 142.360 69.960 143.680 70.250 ;
        RECT 146.030 69.960 147.350 70.250 ;
        RECT 142.360 69.700 142.650 69.960 ;
        RECT 147.060 69.700 147.350 69.960 ;
        RECT 142.360 69.410 147.350 69.700 ;
        RECT 92.560 68.625 93.395 69.135 ;
        RECT 126.760 68.625 127.595 69.135 ;
        RECT 89.265 68.335 93.395 68.625 ;
        RECT 89.265 68.075 89.555 68.335 ;
        RECT 93.105 68.075 93.395 68.335 ;
        RECT 89.265 67.785 90.585 68.075 ;
        RECT 92.075 67.785 93.395 68.075 ;
        RECT 89.265 67.390 89.555 67.785 ;
        RECT 89.925 67.390 90.155 67.595 ;
        RECT 90.355 67.390 90.585 67.595 ;
        RECT 89.265 67.100 90.585 67.390 ;
        RECT 89.265 66.155 89.555 67.100 ;
        RECT 89.925 66.895 90.155 67.100 ;
        RECT 90.355 66.895 90.585 67.100 ;
        RECT 90.770 66.895 91.030 67.595 ;
        RECT 91.200 66.895 91.460 67.595 ;
        RECT 91.630 66.895 91.890 67.595 ;
        RECT 92.075 67.390 92.305 67.595 ;
        RECT 92.505 67.390 92.735 67.595 ;
        RECT 93.105 67.390 93.395 67.785 ;
        RECT 92.075 67.100 93.395 67.390 ;
        RECT 92.075 66.895 92.305 67.100 ;
        RECT 92.505 66.895 92.735 67.100 ;
        RECT 90.230 66.375 91.470 66.705 ;
        RECT 93.105 66.155 93.395 67.100 ;
        RECT 89.265 65.865 93.395 66.155 ;
        RECT 93.895 68.335 98.105 68.625 ;
        RECT 93.895 67.390 94.185 68.335 ;
        RECT 95.885 67.785 97.530 68.115 ;
        RECT 94.595 67.390 94.825 67.595 ;
        RECT 95.025 67.390 95.255 67.595 ;
        RECT 93.895 67.100 95.255 67.390 ;
        RECT 93.895 66.705 94.185 67.100 ;
        RECT 94.595 66.895 94.825 67.100 ;
        RECT 95.025 66.895 95.255 67.100 ;
        RECT 95.440 66.895 95.700 67.595 ;
        RECT 95.870 66.895 96.130 67.595 ;
        RECT 96.300 66.895 96.560 67.595 ;
        RECT 96.745 67.390 96.975 67.595 ;
        RECT 97.175 67.390 97.405 67.595 ;
        RECT 97.815 67.390 98.105 68.335 ;
        RECT 96.745 67.100 98.105 67.390 ;
        RECT 96.745 66.895 96.975 67.100 ;
        RECT 97.175 66.895 97.405 67.100 ;
        RECT 97.815 66.705 98.105 67.100 ;
        RECT 93.895 66.415 95.255 66.705 ;
        RECT 96.745 66.415 98.105 66.705 ;
        RECT 93.895 66.155 94.185 66.415 ;
        RECT 97.815 66.155 98.105 66.415 ;
        RECT 93.895 65.865 98.105 66.155 ;
        RECT 123.465 68.335 127.595 68.625 ;
        RECT 123.465 68.075 123.755 68.335 ;
        RECT 127.305 68.075 127.595 68.335 ;
        RECT 123.465 67.785 124.785 68.075 ;
        RECT 126.275 67.785 127.595 68.075 ;
        RECT 123.465 67.390 123.755 67.785 ;
        RECT 124.125 67.390 124.355 67.595 ;
        RECT 124.555 67.390 124.785 67.595 ;
        RECT 123.465 67.100 124.785 67.390 ;
        RECT 123.465 66.155 123.755 67.100 ;
        RECT 124.125 66.895 124.355 67.100 ;
        RECT 124.555 66.895 124.785 67.100 ;
        RECT 124.970 66.895 125.230 67.595 ;
        RECT 125.400 66.895 125.660 67.595 ;
        RECT 125.830 66.895 126.090 67.595 ;
        RECT 126.275 67.390 126.505 67.595 ;
        RECT 126.705 67.390 126.935 67.595 ;
        RECT 127.305 67.390 127.595 67.785 ;
        RECT 126.275 67.100 127.595 67.390 ;
        RECT 126.275 66.895 126.505 67.100 ;
        RECT 126.705 66.895 126.935 67.100 ;
        RECT 124.430 66.375 125.670 66.705 ;
        RECT 127.305 66.155 127.595 67.100 ;
        RECT 123.465 65.865 127.595 66.155 ;
        RECT 128.095 68.335 132.305 68.625 ;
        RECT 137.070 68.475 139.590 69.410 ;
        RECT 128.095 67.390 128.385 68.335 ;
        RECT 130.085 67.785 131.730 68.115 ;
        RECT 128.795 67.390 129.025 67.595 ;
        RECT 129.225 67.390 129.455 67.595 ;
        RECT 128.095 67.100 129.455 67.390 ;
        RECT 128.095 66.705 128.385 67.100 ;
        RECT 128.795 66.895 129.025 67.100 ;
        RECT 129.225 66.895 129.455 67.100 ;
        RECT 129.640 66.895 129.900 67.595 ;
        RECT 130.070 66.895 130.330 67.595 ;
        RECT 130.500 66.895 130.760 67.595 ;
        RECT 130.945 67.390 131.175 67.595 ;
        RECT 131.375 67.390 131.605 67.595 ;
        RECT 132.015 67.390 132.305 68.335 ;
        RECT 130.945 67.100 132.305 67.390 ;
        RECT 130.945 66.895 131.175 67.100 ;
        RECT 131.375 66.895 131.605 67.100 ;
        RECT 132.015 66.705 132.305 67.100 ;
        RECT 128.095 66.415 129.455 66.705 ;
        RECT 130.945 66.415 132.305 66.705 ;
        RECT 128.095 66.155 128.385 66.415 ;
        RECT 132.015 66.155 132.305 66.415 ;
        RECT 128.095 65.865 132.305 66.155 ;
        RECT 136.790 68.185 147.540 68.475 ;
        RECT 136.790 67.925 137.080 68.185 ;
        RECT 147.250 67.925 147.540 68.185 ;
        RECT 136.790 67.635 139.580 67.925 ;
        RECT 144.750 67.635 147.540 67.925 ;
        RECT 136.790 66.005 137.080 67.635 ;
        RECT 137.475 66.745 137.735 67.445 ;
        RECT 139.755 66.745 140.015 67.445 ;
        RECT 142.035 66.745 142.295 67.445 ;
        RECT 144.315 66.745 144.575 67.445 ;
        RECT 146.595 66.745 146.855 67.445 ;
        RECT 137.960 66.225 144.140 66.555 ;
        RECT 147.250 66.005 147.540 67.635 ;
        RECT 33.520 64.945 38.590 65.235 ;
        RECT 93.895 65.075 96.015 65.865 ;
        RECT 128.095 65.075 130.215 65.865 ;
        RECT 136.790 65.715 147.540 66.005 ;
        RECT 33.520 62.355 33.810 64.945 ;
        RECT 34.220 64.045 34.450 64.545 ;
        RECT 34.650 64.045 34.880 64.545 ;
        RECT 35.080 64.045 35.310 64.545 ;
        RECT 34.205 63.045 34.465 64.045 ;
        RECT 34.635 63.045 34.895 64.045 ;
        RECT 35.065 63.045 35.325 64.045 ;
        RECT 34.220 62.545 34.450 63.045 ;
        RECT 34.650 62.545 34.880 63.045 ;
        RECT 35.080 62.545 35.310 63.045 ;
        RECT 35.495 62.545 35.755 64.545 ;
        RECT 35.940 64.045 36.170 64.545 ;
        RECT 35.925 63.045 36.185 64.045 ;
        RECT 35.940 62.545 36.170 63.045 ;
        RECT 36.355 62.545 36.615 64.545 ;
        RECT 36.800 64.045 37.030 64.545 ;
        RECT 37.230 64.045 37.460 64.545 ;
        RECT 37.660 64.045 37.890 64.545 ;
        RECT 36.785 63.045 37.045 64.045 ;
        RECT 37.215 63.045 37.475 64.045 ;
        RECT 37.645 63.045 37.905 64.045 ;
        RECT 36.800 62.545 37.030 63.045 ;
        RECT 37.230 62.545 37.460 63.045 ;
        RECT 37.660 62.545 37.890 63.045 ;
        RECT 38.300 62.355 38.590 64.945 ;
        RECT 33.520 62.065 35.060 62.355 ;
        RECT 35.330 62.065 36.780 62.355 ;
        RECT 37.050 62.065 38.590 62.355 ;
        RECT 33.520 61.515 33.810 62.065 ;
        RECT 35.890 61.535 36.220 62.065 ;
        RECT 33.520 60.675 33.810 61.225 ;
        RECT 34.215 61.205 36.220 61.535 ;
        RECT 38.300 61.515 38.590 62.065 ;
        RECT 42.670 64.785 144.620 65.075 ;
        RECT 42.670 63.155 42.960 64.785 ;
        RECT 43.355 63.345 43.615 64.045 ;
        RECT 45.635 63.345 45.895 64.045 ;
        RECT 47.915 63.345 48.175 64.045 ;
        RECT 50.185 63.175 50.465 64.045 ;
        RECT 52.475 63.345 52.735 64.045 ;
        RECT 54.745 63.175 55.025 64.045 ;
        RECT 57.035 63.345 57.295 64.045 ;
        RECT 59.305 63.175 59.585 64.045 ;
        RECT 61.595 63.345 61.855 64.045 ;
        RECT 63.865 63.175 64.145 64.045 ;
        RECT 66.155 63.345 66.415 64.045 ;
        RECT 68.425 63.175 68.705 64.045 ;
        RECT 70.715 63.345 70.975 64.045 ;
        RECT 72.995 63.345 73.255 64.045 ;
        RECT 75.275 63.345 75.535 64.045 ;
        RECT 77.555 63.345 77.815 64.045 ;
        RECT 79.835 63.345 80.095 64.045 ;
        RECT 82.115 63.345 82.375 64.045 ;
        RECT 84.395 63.345 84.655 64.045 ;
        RECT 86.675 63.345 86.935 64.045 ;
        RECT 88.955 63.345 89.215 64.045 ;
        RECT 91.235 63.345 91.495 64.045 ;
        RECT 93.515 63.345 93.775 64.045 ;
        RECT 95.795 63.345 96.055 64.045 ;
        RECT 98.075 63.345 98.335 64.045 ;
        RECT 100.355 63.345 100.615 64.045 ;
        RECT 102.635 63.345 102.895 64.045 ;
        RECT 104.915 63.345 105.175 64.045 ;
        RECT 107.195 63.345 107.455 64.045 ;
        RECT 109.475 63.345 109.735 64.045 ;
        RECT 111.755 63.345 112.015 64.045 ;
        RECT 114.035 63.345 114.295 64.045 ;
        RECT 116.315 63.345 116.575 64.045 ;
        RECT 118.595 63.345 118.855 64.045 ;
        RECT 120.875 63.345 121.135 64.045 ;
        RECT 123.155 63.345 123.415 64.045 ;
        RECT 125.435 63.345 125.695 64.045 ;
        RECT 127.715 63.345 127.975 64.045 ;
        RECT 129.995 63.345 130.255 64.045 ;
        RECT 132.275 63.345 132.535 64.045 ;
        RECT 134.555 63.345 134.815 64.045 ;
        RECT 136.835 63.345 137.095 64.045 ;
        RECT 139.115 63.345 139.375 64.045 ;
        RECT 141.395 63.345 141.655 64.045 ;
        RECT 143.675 63.345 143.935 64.045 ;
        RECT 42.670 62.865 47.740 63.155 ;
        RECT 42.670 61.785 42.960 62.865 ;
        RECT 48.350 62.845 138.940 63.175 ;
        RECT 144.330 63.155 144.620 64.785 ;
        RECT 139.550 62.865 144.620 63.155 ;
        RECT 43.355 61.975 43.615 62.675 ;
        RECT 45.635 61.975 45.895 62.675 ;
        RECT 47.915 61.975 48.175 62.675 ;
        RECT 50.185 61.805 50.465 62.845 ;
        RECT 52.475 61.975 52.735 62.675 ;
        RECT 54.745 61.805 55.025 62.845 ;
        RECT 57.035 61.975 57.295 62.675 ;
        RECT 59.305 61.805 59.585 62.845 ;
        RECT 61.595 61.975 61.855 62.675 ;
        RECT 63.865 61.805 64.145 62.845 ;
        RECT 66.155 61.975 66.415 62.675 ;
        RECT 68.425 61.805 68.705 62.845 ;
        RECT 70.715 61.975 70.975 62.675 ;
        RECT 72.995 61.975 73.255 62.675 ;
        RECT 75.275 61.975 75.535 62.675 ;
        RECT 77.555 61.975 77.815 62.675 ;
        RECT 79.835 61.975 80.095 62.675 ;
        RECT 82.115 61.975 82.375 62.675 ;
        RECT 84.395 61.975 84.655 62.675 ;
        RECT 86.675 61.975 86.935 62.675 ;
        RECT 88.955 61.975 89.215 62.675 ;
        RECT 91.235 61.975 91.495 62.675 ;
        RECT 93.515 61.975 93.775 62.675 ;
        RECT 95.795 61.975 96.055 62.675 ;
        RECT 98.075 61.975 98.335 62.675 ;
        RECT 100.355 61.975 100.615 62.675 ;
        RECT 102.635 61.975 102.895 62.675 ;
        RECT 104.915 61.975 105.175 62.675 ;
        RECT 107.195 61.975 107.455 62.675 ;
        RECT 109.475 61.975 109.735 62.675 ;
        RECT 111.755 61.975 112.015 62.675 ;
        RECT 114.035 61.975 114.295 62.675 ;
        RECT 116.315 61.975 116.575 62.675 ;
        RECT 118.595 61.975 118.855 62.675 ;
        RECT 120.875 61.975 121.135 62.675 ;
        RECT 123.155 61.975 123.415 62.675 ;
        RECT 125.435 61.975 125.695 62.675 ;
        RECT 127.715 61.975 127.975 62.675 ;
        RECT 129.995 61.975 130.255 62.675 ;
        RECT 132.275 61.975 132.535 62.675 ;
        RECT 134.555 61.975 134.815 62.675 ;
        RECT 136.835 61.975 137.095 62.675 ;
        RECT 139.115 61.975 139.375 62.675 ;
        RECT 141.395 61.975 141.655 62.675 ;
        RECT 143.675 61.975 143.935 62.675 ;
        RECT 42.670 61.495 47.740 61.785 ;
        RECT 35.890 60.675 36.220 61.205 ;
        RECT 38.300 60.675 38.590 61.225 ;
        RECT 33.520 60.385 35.060 60.675 ;
        RECT 35.330 60.385 36.780 60.675 ;
        RECT 37.050 60.385 38.590 60.675 ;
        RECT 33.520 58.820 33.810 60.385 ;
        RECT 34.205 59.195 34.465 60.195 ;
        RECT 34.635 59.195 34.895 60.195 ;
        RECT 35.065 59.195 35.325 60.195 ;
        RECT 35.495 59.195 35.755 60.195 ;
        RECT 35.925 59.195 36.185 60.195 ;
        RECT 36.355 59.195 36.615 60.195 ;
        RECT 36.785 59.195 37.045 60.195 ;
        RECT 37.215 59.195 37.475 60.195 ;
        RECT 37.645 59.195 37.905 60.195 ;
        RECT 38.300 58.820 38.590 60.385 ;
        RECT 42.670 59.865 42.960 61.495 ;
        RECT 48.350 61.475 138.940 61.805 ;
        RECT 144.330 61.785 144.620 62.865 ;
        RECT 139.550 61.495 144.620 61.785 ;
        RECT 43.355 60.605 43.615 61.305 ;
        RECT 45.635 60.605 45.895 61.305 ;
        RECT 47.915 60.605 48.175 61.305 ;
        RECT 50.185 60.605 50.465 61.475 ;
        RECT 52.475 60.605 52.735 61.305 ;
        RECT 54.745 60.605 55.025 61.475 ;
        RECT 57.035 60.605 57.295 61.305 ;
        RECT 59.305 60.605 59.585 61.475 ;
        RECT 61.595 60.605 61.855 61.305 ;
        RECT 63.865 60.605 64.145 61.475 ;
        RECT 66.155 60.605 66.415 61.305 ;
        RECT 68.425 60.605 68.705 61.475 ;
        RECT 70.715 60.605 70.975 61.305 ;
        RECT 72.995 60.605 73.255 61.305 ;
        RECT 75.275 60.605 75.535 61.305 ;
        RECT 77.555 60.605 77.815 61.305 ;
        RECT 79.835 60.605 80.095 61.305 ;
        RECT 82.115 60.605 82.375 61.305 ;
        RECT 84.395 60.605 84.655 61.305 ;
        RECT 86.675 60.605 86.935 61.305 ;
        RECT 88.955 60.605 89.215 61.305 ;
        RECT 91.235 60.605 91.495 61.305 ;
        RECT 93.515 60.605 93.775 61.305 ;
        RECT 95.795 60.605 96.055 61.305 ;
        RECT 98.075 60.605 98.335 61.305 ;
        RECT 100.355 60.605 100.615 61.305 ;
        RECT 102.635 60.605 102.895 61.305 ;
        RECT 104.915 60.605 105.175 61.305 ;
        RECT 107.195 60.605 107.455 61.305 ;
        RECT 109.475 60.605 109.735 61.305 ;
        RECT 111.755 60.605 112.015 61.305 ;
        RECT 114.035 60.605 114.295 61.305 ;
        RECT 116.315 60.605 116.575 61.305 ;
        RECT 118.595 60.605 118.855 61.305 ;
        RECT 120.875 60.605 121.135 61.305 ;
        RECT 123.155 60.605 123.415 61.305 ;
        RECT 125.435 60.605 125.695 61.305 ;
        RECT 127.715 60.605 127.975 61.305 ;
        RECT 129.995 60.605 130.255 61.305 ;
        RECT 132.275 60.605 132.535 61.305 ;
        RECT 134.555 60.605 134.815 61.305 ;
        RECT 136.835 60.605 137.095 61.305 ;
        RECT 139.115 60.605 139.375 61.305 ;
        RECT 141.395 60.605 141.655 61.305 ;
        RECT 143.675 60.605 143.935 61.305 ;
        RECT 144.330 59.865 144.620 61.495 ;
        RECT 42.670 59.575 144.620 59.865 ;
        RECT 33.520 58.530 38.590 58.820 ;
        RECT 55.920 53.380 95.710 53.670 ;
        RECT 55.920 51.450 56.210 53.380 ;
        RECT 77.680 52.830 81.630 53.160 ;
        RECT 65.845 51.640 66.105 52.640 ;
        RECT 68.125 51.640 68.385 52.640 ;
        RECT 70.405 51.640 70.665 52.640 ;
        RECT 72.685 51.640 72.945 52.640 ;
        RECT 74.965 51.640 75.225 52.640 ;
        RECT 77.245 51.640 77.505 52.640 ;
        RECT 79.525 51.640 79.785 52.640 ;
        RECT 81.805 51.640 82.065 52.640 ;
        RECT 84.085 51.640 84.345 52.640 ;
        RECT 86.365 51.640 86.625 52.640 ;
        RECT 88.645 51.640 88.905 52.640 ;
        RECT 90.925 51.640 91.185 52.640 ;
        RECT 93.205 51.640 93.465 52.640 ;
        RECT 95.420 51.450 95.710 53.380 ;
        RECT 55.920 51.160 77.070 51.450 ;
        RECT 82.240 51.160 95.710 51.450 ;
        RECT 55.920 49.530 56.210 51.160 ;
        RECT 95.420 49.530 95.710 51.160 ;
        RECT 55.920 49.240 57.990 49.530 ;
        RECT 63.160 49.240 65.670 49.530 ;
        RECT 66.280 49.240 67.950 49.530 ;
        RECT 68.560 49.240 70.230 49.530 ;
        RECT 70.840 49.240 72.510 49.530 ;
        RECT 73.120 49.240 74.790 49.530 ;
        RECT 75.400 49.240 77.070 49.530 ;
        RECT 77.680 49.240 79.350 49.530 ;
        RECT 79.960 49.240 81.630 49.530 ;
        RECT 82.240 49.240 83.910 49.530 ;
        RECT 84.520 49.240 86.190 49.530 ;
        RECT 86.800 49.240 88.470 49.530 ;
        RECT 89.080 49.240 90.750 49.530 ;
        RECT 91.360 49.240 93.030 49.530 ;
        RECT 93.640 49.240 95.710 49.530 ;
        RECT 55.920 47.310 56.210 49.240 ;
        RECT 56.605 48.050 56.865 49.050 ;
        RECT 57.385 48.050 57.645 49.050 ;
        RECT 58.165 48.050 58.425 49.050 ;
        RECT 60.445 48.050 60.705 49.050 ;
        RECT 62.725 48.050 62.985 49.050 ;
        RECT 63.490 48.050 63.780 49.240 ;
        RECT 64.270 48.050 64.560 49.240 ;
        RECT 65.050 48.050 65.340 49.240 ;
        RECT 65.845 48.050 66.105 49.050 ;
        RECT 68.125 48.050 68.385 49.050 ;
        RECT 70.405 48.050 70.665 49.050 ;
        RECT 72.685 48.050 72.945 49.050 ;
        RECT 74.965 48.050 75.225 49.050 ;
        RECT 77.245 48.050 77.505 49.050 ;
        RECT 79.525 48.050 79.785 49.050 ;
        RECT 81.805 48.050 82.065 49.050 ;
        RECT 84.085 48.050 84.345 49.050 ;
        RECT 86.365 48.050 86.625 49.050 ;
        RECT 88.645 48.050 88.905 49.050 ;
        RECT 90.925 48.050 91.185 49.050 ;
        RECT 93.205 48.050 93.465 49.050 ;
        RECT 93.985 48.050 94.245 49.050 ;
        RECT 94.765 48.050 95.025 49.050 ;
        RECT 58.600 47.530 62.550 47.860 ;
        RECT 66.280 47.530 79.350 47.860 ;
        RECT 79.960 47.530 93.030 47.860 ;
        RECT 95.420 47.310 95.710 49.240 ;
        RECT 55.920 47.020 95.710 47.310 ;
        RECT 94.080 45.875 118.510 46.165 ;
        RECT 55.920 45.125 65.230 45.415 ;
        RECT 55.920 43.695 56.210 45.125 ;
        RECT 58.600 44.575 62.550 44.905 ;
        RECT 56.605 43.885 56.865 44.385 ;
        RECT 57.385 43.885 57.645 44.385 ;
        RECT 58.165 43.885 58.425 44.385 ;
        RECT 60.445 43.885 60.705 44.385 ;
        RECT 62.725 43.885 62.985 44.385 ;
        RECT 63.505 43.885 63.765 44.385 ;
        RECT 64.285 43.885 64.545 44.385 ;
        RECT 64.940 43.695 65.230 45.125 ;
        RECT 55.920 43.405 57.990 43.695 ;
        RECT 63.160 43.405 65.230 43.695 ;
        RECT 55.920 43.145 56.210 43.405 ;
        RECT 64.940 43.145 65.230 43.405 ;
        RECT 55.920 42.855 65.230 43.145 ;
        RECT 69.130 45.125 90.120 45.415 ;
        RECT 69.130 44.865 69.420 45.125 ;
        RECT 69.130 44.575 72.245 44.865 ;
        RECT 72.675 44.575 76.760 44.905 ;
        RECT 77.335 44.575 81.925 44.865 ;
        RECT 82.490 44.580 86.440 44.910 ;
        RECT 89.830 44.865 90.120 45.125 ;
        RECT 82.490 44.575 84.160 44.580 ;
        RECT 84.770 44.575 86.440 44.580 ;
        RECT 87.015 44.575 90.120 44.865 ;
        RECT 69.130 43.715 69.420 44.575 ;
        RECT 69.815 43.885 70.075 44.385 ;
        RECT 71.095 43.885 71.355 44.385 ;
        RECT 72.375 43.885 72.635 44.385 ;
        RECT 69.130 43.425 72.245 43.715 ;
        RECT 74.635 43.695 74.925 44.575 ;
        RECT 76.935 43.885 77.195 44.385 ;
        RECT 78.205 43.715 78.485 44.575 ;
        RECT 79.485 43.715 79.765 44.575 ;
        RECT 80.765 43.715 81.045 44.575 ;
        RECT 82.055 43.885 82.315 44.385 ;
        RECT 84.335 43.885 84.595 44.385 ;
        RECT 86.615 43.885 86.875 44.385 ;
        RECT 87.895 43.885 88.155 44.385 ;
        RECT 89.175 43.885 89.435 44.385 ;
        RECT 89.830 43.715 90.120 44.575 ;
        RECT 69.130 43.145 69.420 43.425 ;
        RECT 70.215 43.405 72.245 43.425 ;
        RECT 72.810 43.365 76.760 43.695 ;
        RECT 77.335 43.425 81.925 43.715 ;
        RECT 77.335 43.405 79.365 43.425 ;
        RECT 79.895 43.405 81.925 43.425 ;
        RECT 87.015 43.425 90.120 43.715 ;
        RECT 87.015 43.405 89.045 43.425 ;
        RECT 89.830 43.145 90.120 43.425 ;
        RECT 69.130 42.855 90.120 43.145 ;
        RECT 94.080 44.285 94.370 45.875 ;
        RECT 94.765 44.475 95.025 45.475 ;
        RECT 97.045 44.475 97.305 45.475 ;
        RECT 99.325 44.475 99.585 45.475 ;
        RECT 101.605 44.475 101.865 45.475 ;
        RECT 103.885 44.475 104.145 45.475 ;
        RECT 106.165 44.475 106.425 45.475 ;
        RECT 108.445 44.475 108.705 45.475 ;
        RECT 110.725 44.475 110.985 45.475 ;
        RECT 113.005 44.475 113.265 45.475 ;
        RECT 115.285 44.475 115.545 45.475 ;
        RECT 117.565 44.475 117.825 45.475 ;
        RECT 118.220 44.285 118.510 45.875 ;
        RECT 94.080 43.995 99.150 44.285 ;
        RECT 94.080 42.445 94.370 43.995 ;
        RECT 99.760 43.955 103.710 44.285 ;
        RECT 104.320 43.955 108.270 44.285 ;
        RECT 108.880 43.955 112.830 44.285 ;
        RECT 113.440 43.995 118.510 44.285 ;
        RECT 101.595 42.450 101.875 42.765 ;
        RECT 104.320 42.450 104.650 43.955 ;
        RECT 69.130 41.370 90.120 41.660 ;
        RECT 69.130 41.090 69.420 41.370 ;
        RECT 70.215 41.090 72.245 41.110 ;
        RECT 69.130 40.800 72.245 41.090 ;
        RECT 72.810 40.820 76.760 41.150 ;
        RECT 77.335 41.090 79.365 41.110 ;
        RECT 79.895 41.090 81.925 41.110 ;
        RECT 77.335 40.800 81.925 41.090 ;
        RECT 87.015 41.090 89.045 41.110 ;
        RECT 89.830 41.090 90.120 41.370 ;
        RECT 87.015 40.800 90.120 41.090 ;
        RECT 69.130 39.460 69.420 40.800 ;
        RECT 69.815 39.630 70.075 40.630 ;
        RECT 71.095 39.630 71.355 40.630 ;
        RECT 72.375 39.630 72.635 40.630 ;
        RECT 74.670 39.460 74.935 40.630 ;
        RECT 76.935 39.630 77.195 40.630 ;
        RECT 78.205 39.460 78.485 40.800 ;
        RECT 79.485 39.460 79.765 40.800 ;
        RECT 80.765 39.460 81.045 40.800 ;
        RECT 82.055 39.630 82.315 40.630 ;
        RECT 84.350 39.460 84.625 40.630 ;
        RECT 86.615 39.630 86.875 40.630 ;
        RECT 87.895 39.630 88.155 40.630 ;
        RECT 89.175 39.630 89.435 40.630 ;
        RECT 89.830 39.460 90.120 40.800 ;
        RECT 94.080 41.155 94.370 42.180 ;
        RECT 101.595 42.120 104.650 42.450 ;
        RECT 101.595 41.805 101.875 42.120 ;
        RECT 104.320 41.195 104.650 42.120 ;
        RECT 106.155 42.450 106.435 42.765 ;
        RECT 108.880 42.450 109.210 43.955 ;
        RECT 106.155 42.120 109.210 42.450 ;
        RECT 118.220 42.445 118.510 43.995 ;
        RECT 124.400 45.860 129.470 46.150 ;
        RECT 124.400 43.270 124.690 45.860 ;
        RECT 125.100 44.960 125.330 45.460 ;
        RECT 125.530 44.960 125.760 45.460 ;
        RECT 125.960 44.960 126.190 45.460 ;
        RECT 125.085 43.960 125.345 44.960 ;
        RECT 125.515 43.960 125.775 44.960 ;
        RECT 125.945 43.960 126.205 44.960 ;
        RECT 125.100 43.460 125.330 43.960 ;
        RECT 125.530 43.460 125.760 43.960 ;
        RECT 125.960 43.460 126.190 43.960 ;
        RECT 126.375 43.460 126.635 45.460 ;
        RECT 126.820 44.960 127.050 45.460 ;
        RECT 126.805 43.960 127.065 44.960 ;
        RECT 126.820 43.460 127.050 43.960 ;
        RECT 127.235 43.460 127.495 45.460 ;
        RECT 127.680 44.960 127.910 45.460 ;
        RECT 128.110 44.960 128.340 45.460 ;
        RECT 128.540 44.960 128.770 45.460 ;
        RECT 127.665 43.960 127.925 44.960 ;
        RECT 128.095 43.960 128.355 44.960 ;
        RECT 128.525 43.960 128.785 44.960 ;
        RECT 127.680 43.460 127.910 43.960 ;
        RECT 128.110 43.460 128.340 43.960 ;
        RECT 128.540 43.460 128.770 43.960 ;
        RECT 129.180 43.270 129.470 45.860 ;
        RECT 124.400 42.980 125.940 43.270 ;
        RECT 126.210 42.980 127.660 43.270 ;
        RECT 127.930 42.980 129.470 43.270 ;
        RECT 124.400 42.430 124.690 42.980 ;
        RECT 126.770 42.450 127.100 42.980 ;
        RECT 106.155 41.805 106.435 42.120 ;
        RECT 108.880 41.195 109.210 42.120 ;
        RECT 94.080 40.865 99.150 41.155 ;
        RECT 99.760 40.865 103.710 41.195 ;
        RECT 104.320 40.865 108.270 41.195 ;
        RECT 108.880 40.865 112.830 41.195 ;
        RECT 118.220 41.155 118.510 42.180 ;
        RECT 113.440 40.865 118.510 41.155 ;
        RECT 94.080 39.775 94.370 40.865 ;
        RECT 94.765 40.175 95.025 40.675 ;
        RECT 97.045 40.175 97.305 40.675 ;
        RECT 99.325 40.175 99.585 40.675 ;
        RECT 101.605 40.175 101.865 40.675 ;
        RECT 103.885 40.175 104.145 40.675 ;
        RECT 106.165 40.175 106.425 40.675 ;
        RECT 108.445 40.175 108.705 40.675 ;
        RECT 110.725 40.175 110.985 40.675 ;
        RECT 113.005 40.175 113.265 40.675 ;
        RECT 115.285 40.175 115.545 40.675 ;
        RECT 117.565 40.175 117.825 40.675 ;
        RECT 118.220 39.775 118.510 40.865 ;
        RECT 94.080 39.485 118.510 39.775 ;
        RECT 124.400 41.590 124.690 42.140 ;
        RECT 125.095 42.120 127.100 42.450 ;
        RECT 129.180 42.430 129.470 42.980 ;
        RECT 135.060 45.860 144.430 46.150 ;
        RECT 135.060 43.270 135.350 45.860 ;
        RECT 135.760 44.960 135.990 45.460 ;
        RECT 136.190 44.960 136.420 45.460 ;
        RECT 136.620 44.960 136.850 45.460 ;
        RECT 135.745 43.960 136.005 44.960 ;
        RECT 136.175 43.960 136.435 44.960 ;
        RECT 136.605 43.960 136.865 44.960 ;
        RECT 135.760 43.460 135.990 43.960 ;
        RECT 136.190 43.460 136.420 43.960 ;
        RECT 136.620 43.460 136.850 43.960 ;
        RECT 137.035 43.460 137.295 45.460 ;
        RECT 137.480 44.960 137.710 45.460 ;
        RECT 137.465 43.960 137.725 44.960 ;
        RECT 137.480 43.460 137.710 43.960 ;
        RECT 137.895 43.460 138.155 45.460 ;
        RECT 138.340 44.960 138.570 45.460 ;
        RECT 138.325 43.960 138.585 44.960 ;
        RECT 138.340 43.460 138.570 43.960 ;
        RECT 138.755 43.460 139.015 45.460 ;
        RECT 139.200 44.960 139.430 45.460 ;
        RECT 139.185 43.960 139.445 44.960 ;
        RECT 139.200 43.460 139.430 43.960 ;
        RECT 139.615 43.460 139.875 45.460 ;
        RECT 140.060 44.960 140.290 45.460 ;
        RECT 140.045 43.960 140.305 44.960 ;
        RECT 140.060 43.460 140.290 43.960 ;
        RECT 140.475 43.460 140.735 45.460 ;
        RECT 140.920 44.960 141.150 45.460 ;
        RECT 140.905 43.960 141.165 44.960 ;
        RECT 140.920 43.460 141.150 43.960 ;
        RECT 141.335 43.460 141.595 45.460 ;
        RECT 141.780 44.960 142.010 45.460 ;
        RECT 141.765 43.960 142.025 44.960 ;
        RECT 141.780 43.460 142.010 43.960 ;
        RECT 142.195 43.460 142.455 45.460 ;
        RECT 142.640 44.960 142.870 45.460 ;
        RECT 143.070 44.960 143.300 45.460 ;
        RECT 143.500 44.960 143.730 45.460 ;
        RECT 142.625 43.960 142.885 44.960 ;
        RECT 143.055 43.960 143.315 44.960 ;
        RECT 143.485 43.960 143.745 44.960 ;
        RECT 142.640 43.460 142.870 43.960 ;
        RECT 143.070 43.460 143.300 43.960 ;
        RECT 143.500 43.460 143.730 43.960 ;
        RECT 144.140 43.270 144.430 45.860 ;
        RECT 135.060 42.980 136.600 43.270 ;
        RECT 136.870 42.980 138.320 43.270 ;
        RECT 138.590 42.980 142.620 43.270 ;
        RECT 142.890 42.980 144.430 43.270 ;
        RECT 135.060 42.430 135.350 42.980 ;
        RECT 137.415 42.450 137.745 42.980 ;
        RECT 126.770 41.590 127.100 42.120 ;
        RECT 129.180 41.590 129.470 42.140 ;
        RECT 124.400 41.300 125.940 41.590 ;
        RECT 126.210 41.300 127.660 41.590 ;
        RECT 127.930 41.300 129.470 41.590 ;
        RECT 124.400 39.735 124.690 41.300 ;
        RECT 125.085 40.110 125.345 41.110 ;
        RECT 125.515 40.110 125.775 41.110 ;
        RECT 125.945 40.110 126.205 41.110 ;
        RECT 126.375 40.110 126.635 41.110 ;
        RECT 126.805 40.110 127.065 41.110 ;
        RECT 127.235 40.110 127.495 41.110 ;
        RECT 127.665 40.110 127.925 41.110 ;
        RECT 128.095 40.110 128.355 41.110 ;
        RECT 128.525 40.110 128.785 41.110 ;
        RECT 129.180 39.735 129.470 41.300 ;
        RECT 69.130 39.170 72.245 39.460 ;
        RECT 69.130 38.890 69.420 39.170 ;
        RECT 70.215 39.150 72.245 39.170 ;
        RECT 72.810 39.130 76.760 39.460 ;
        RECT 77.335 39.170 81.925 39.460 ;
        RECT 77.335 39.150 79.365 39.170 ;
        RECT 79.895 39.150 81.925 39.170 ;
        RECT 82.490 39.130 86.440 39.460 ;
        RECT 87.015 39.170 90.120 39.460 ;
        RECT 124.400 39.445 129.470 39.735 ;
        RECT 135.060 41.590 135.350 42.140 ;
        RECT 135.755 42.120 137.745 42.450 ;
        RECT 137.415 41.590 137.745 42.120 ;
        RECT 137.885 42.450 138.165 42.765 ;
        RECT 140.440 42.450 140.770 42.980 ;
        RECT 137.885 42.120 140.770 42.450 ;
        RECT 144.140 42.430 144.430 42.980 ;
        RECT 137.885 41.805 138.165 42.120 ;
        RECT 140.440 41.590 140.770 42.120 ;
        RECT 144.140 41.590 144.430 42.140 ;
        RECT 135.060 41.300 136.600 41.590 ;
        RECT 136.870 41.300 138.320 41.590 ;
        RECT 138.590 41.300 142.620 41.590 ;
        RECT 142.890 41.300 144.430 41.590 ;
        RECT 135.060 39.735 135.350 41.300 ;
        RECT 135.745 40.110 136.005 41.110 ;
        RECT 136.175 40.110 136.435 41.110 ;
        RECT 136.605 40.110 136.865 41.110 ;
        RECT 137.035 40.110 137.295 41.110 ;
        RECT 137.465 40.110 137.725 41.110 ;
        RECT 137.895 40.110 138.155 41.110 ;
        RECT 138.325 40.110 138.585 41.110 ;
        RECT 138.755 40.110 139.015 41.110 ;
        RECT 139.185 40.110 139.445 41.110 ;
        RECT 139.615 40.110 139.875 41.110 ;
        RECT 140.045 40.110 140.305 41.110 ;
        RECT 140.475 40.110 140.735 41.110 ;
        RECT 140.905 40.110 141.165 41.110 ;
        RECT 141.335 40.110 141.595 41.110 ;
        RECT 141.765 40.110 142.025 41.110 ;
        RECT 142.195 40.110 142.455 41.110 ;
        RECT 142.625 40.110 142.885 41.110 ;
        RECT 143.055 40.110 143.315 41.110 ;
        RECT 143.485 40.110 143.745 41.110 ;
        RECT 144.140 39.735 144.430 41.300 ;
        RECT 135.060 39.445 144.430 39.735 ;
        RECT 87.015 39.150 89.045 39.170 ;
        RECT 89.830 38.890 90.120 39.170 ;
        RECT 69.130 38.600 90.120 38.890 ;
        RECT 124.750 37.855 129.820 38.145 ;
        RECT 64.640 36.970 94.670 37.260 ;
        RECT 64.640 35.540 64.930 36.970 ;
        RECT 66.280 36.420 76.790 36.750 ;
        RECT 77.365 36.420 81.955 36.710 ;
        RECT 82.520 36.420 93.030 36.750 ;
        RECT 65.285 35.730 65.545 36.230 ;
        RECT 66.580 35.540 66.810 36.230 ;
        RECT 67.845 35.730 68.105 36.230 ;
        RECT 70.125 35.730 70.385 36.230 ;
        RECT 72.405 35.730 72.665 36.230 ;
        RECT 74.685 35.730 74.945 36.230 ;
        RECT 76.965 35.730 77.225 36.230 ;
        RECT 78.235 35.540 78.515 36.420 ;
        RECT 79.515 35.540 79.795 36.420 ;
        RECT 80.795 35.540 81.075 36.420 ;
        RECT 82.085 35.730 82.345 36.230 ;
        RECT 84.365 35.730 84.625 36.230 ;
        RECT 86.645 35.730 86.905 36.230 ;
        RECT 88.925 35.730 89.185 36.230 ;
        RECT 91.205 35.730 91.465 36.230 ;
        RECT 92.500 35.540 92.730 36.230 ;
        RECT 93.765 35.730 94.025 36.230 ;
        RECT 94.380 35.540 94.670 36.970 ;
        RECT 64.640 35.250 67.715 35.540 ;
        RECT 68.280 35.250 69.950 35.540 ;
        RECT 70.560 35.250 72.230 35.540 ;
        RECT 72.840 35.250 74.510 35.540 ;
        RECT 75.120 35.250 76.790 35.540 ;
        RECT 77.365 35.250 81.955 35.540 ;
        RECT 82.520 35.250 84.190 35.540 ;
        RECT 84.800 35.250 86.470 35.540 ;
        RECT 87.080 35.250 88.750 35.540 ;
        RECT 89.360 35.250 91.030 35.540 ;
        RECT 91.605 35.250 94.670 35.540 ;
        RECT 64.640 33.970 64.930 35.250 ;
        RECT 94.380 33.970 94.670 35.250 ;
        RECT 124.750 35.925 125.040 37.855 ;
        RECT 125.700 37.305 126.290 37.595 ;
        RECT 126.560 37.305 127.150 37.635 ;
        RECT 127.420 37.305 128.010 37.595 ;
        RECT 128.280 37.305 128.870 37.595 ;
        RECT 125.450 36.965 125.680 37.115 ;
        RECT 125.880 36.965 126.110 37.115 ;
        RECT 126.310 36.965 126.540 37.115 ;
        RECT 125.435 36.115 125.695 36.965 ;
        RECT 125.865 36.115 126.125 36.965 ;
        RECT 126.295 36.115 126.555 36.965 ;
        RECT 126.725 36.115 126.985 37.115 ;
        RECT 127.170 36.965 127.400 37.115 ;
        RECT 127.155 36.115 127.415 36.965 ;
        RECT 127.585 36.115 127.845 37.115 ;
        RECT 128.030 36.965 128.260 37.115 ;
        RECT 128.460 36.965 128.690 37.115 ;
        RECT 128.890 36.965 129.120 37.115 ;
        RECT 129.530 36.965 129.820 37.855 ;
        RECT 128.015 36.115 128.275 36.965 ;
        RECT 128.445 36.115 128.705 36.965 ;
        RECT 128.875 36.115 129.135 36.965 ;
        RECT 129.525 36.115 129.820 36.965 ;
        RECT 129.530 35.925 129.820 36.115 ;
        RECT 124.750 35.635 126.290 35.925 ;
        RECT 126.560 35.635 127.150 35.925 ;
        RECT 127.420 35.635 128.010 35.925 ;
        RECT 128.280 35.635 129.820 35.925 ;
        RECT 124.750 35.170 125.040 35.635 ;
        RECT 127.550 35.130 127.880 35.635 ;
        RECT 129.530 35.170 129.820 35.635 ;
        RECT 135.060 37.515 144.430 37.805 ;
        RECT 135.060 35.950 135.350 37.515 ;
        RECT 135.745 36.140 136.005 37.140 ;
        RECT 136.175 36.140 136.435 37.140 ;
        RECT 136.605 36.140 136.865 37.140 ;
        RECT 137.035 36.140 137.295 37.140 ;
        RECT 137.465 36.140 137.725 37.140 ;
        RECT 137.895 36.140 138.155 37.140 ;
        RECT 138.325 36.140 138.585 37.140 ;
        RECT 138.755 36.140 139.015 37.140 ;
        RECT 139.185 36.140 139.445 37.140 ;
        RECT 139.615 36.140 139.875 37.140 ;
        RECT 140.045 36.140 140.305 37.140 ;
        RECT 140.475 36.140 140.735 37.140 ;
        RECT 140.905 36.140 141.165 37.140 ;
        RECT 141.335 36.140 141.595 37.140 ;
        RECT 141.765 36.140 142.025 37.140 ;
        RECT 142.195 36.140 142.455 37.140 ;
        RECT 142.625 36.140 142.885 37.140 ;
        RECT 143.055 36.140 143.315 37.140 ;
        RECT 143.485 36.140 143.745 37.140 ;
        RECT 144.140 35.950 144.430 37.515 ;
        RECT 135.060 35.660 136.600 35.950 ;
        RECT 136.870 35.660 138.320 35.950 ;
        RECT 138.590 35.660 142.620 35.950 ;
        RECT 142.890 35.660 144.430 35.950 ;
        RECT 125.505 34.800 127.880 35.130 ;
        RECT 135.060 35.110 135.350 35.660 ;
        RECT 137.415 35.130 137.745 35.660 ;
        RECT 64.640 33.680 72.115 33.970 ;
        RECT 87.205 33.680 94.670 33.970 ;
        RECT 64.640 32.800 64.930 33.680 ;
        RECT 65.685 32.990 65.945 33.490 ;
        RECT 68.965 32.990 69.225 33.490 ;
        RECT 72.245 32.990 72.505 33.490 ;
        RECT 79.525 32.990 79.785 33.490 ;
        RECT 86.805 32.990 87.065 33.490 ;
        RECT 90.085 32.990 90.345 33.490 ;
        RECT 93.365 32.990 93.625 33.490 ;
        RECT 94.380 32.800 94.670 33.680 ;
        RECT 64.640 32.510 72.115 32.800 ;
        RECT 64.640 32.250 64.930 32.510 ;
        RECT 72.660 32.470 86.650 32.800 ;
        RECT 87.205 32.510 94.670 32.800 ;
        RECT 94.380 32.250 94.670 32.510 ;
        RECT 64.640 31.960 94.670 32.250 ;
        RECT 124.750 34.295 125.040 34.760 ;
        RECT 127.550 34.335 127.880 34.800 ;
        RECT 124.750 34.005 126.290 34.295 ;
        RECT 126.560 34.005 128.010 34.335 ;
        RECT 129.530 34.295 129.820 34.760 ;
        RECT 128.280 34.005 129.820 34.295 ;
        RECT 124.750 30.935 125.040 34.005 ;
        RECT 125.450 33.740 125.680 33.815 ;
        RECT 125.880 33.740 126.110 33.815 ;
        RECT 125.435 32.890 125.695 33.740 ;
        RECT 125.865 32.890 126.125 33.740 ;
        RECT 125.450 32.815 125.680 32.890 ;
        RECT 125.880 32.815 126.110 32.890 ;
        RECT 126.295 32.815 126.555 33.815 ;
        RECT 126.725 32.815 126.985 33.815 ;
        RECT 127.155 32.815 127.415 33.815 ;
        RECT 127.585 32.815 127.845 33.815 ;
        RECT 128.015 32.815 128.275 33.815 ;
        RECT 128.460 33.740 128.690 33.815 ;
        RECT 128.890 33.740 129.120 33.815 ;
        RECT 129.530 33.740 129.820 34.005 ;
        RECT 128.445 32.890 128.705 33.740 ;
        RECT 128.875 32.890 129.135 33.740 ;
        RECT 129.525 32.890 129.820 33.740 ;
        RECT 128.460 32.815 128.690 32.890 ;
        RECT 128.890 32.815 129.120 32.890 ;
        RECT 129.530 32.165 129.820 32.890 ;
        RECT 125.435 31.315 125.695 32.165 ;
        RECT 125.865 31.315 126.125 32.165 ;
        RECT 126.295 31.315 126.555 32.165 ;
        RECT 125.450 31.165 125.680 31.315 ;
        RECT 125.880 31.165 126.110 31.315 ;
        RECT 126.310 31.165 126.540 31.315 ;
        RECT 126.725 31.165 126.985 32.165 ;
        RECT 127.155 31.315 127.415 32.165 ;
        RECT 127.170 31.165 127.400 31.315 ;
        RECT 127.585 31.165 127.845 32.165 ;
        RECT 128.015 31.315 128.275 32.165 ;
        RECT 128.445 31.315 128.705 32.165 ;
        RECT 128.875 31.315 129.135 32.165 ;
        RECT 129.525 31.315 129.820 32.165 ;
        RECT 128.030 31.165 128.260 31.315 ;
        RECT 128.460 31.165 128.690 31.315 ;
        RECT 128.890 31.165 129.120 31.315 ;
        RECT 125.700 30.935 126.290 30.975 ;
        RECT 124.750 30.645 126.290 30.935 ;
        RECT 126.560 30.645 128.010 30.975 ;
        RECT 128.280 30.935 128.870 30.975 ;
        RECT 129.530 30.935 129.820 31.315 ;
        RECT 128.280 30.645 129.820 30.935 ;
        RECT 124.750 30.425 125.040 30.645 ;
        RECT 129.530 30.425 129.820 30.645 ;
        RECT 124.750 30.135 129.820 30.425 ;
        RECT 124.750 29.915 125.040 30.135 ;
        RECT 129.530 29.915 129.820 30.135 ;
        RECT 124.750 29.625 126.290 29.915 ;
        RECT 64.640 28.540 94.670 28.830 ;
        RECT 64.640 28.280 64.930 28.540 ;
        RECT 64.640 27.990 72.115 28.280 ;
        RECT 72.660 27.990 86.650 28.320 ;
        RECT 94.380 28.280 94.670 28.540 ;
        RECT 87.205 27.990 94.670 28.280 ;
        RECT 64.640 27.110 64.930 27.990 ;
        RECT 65.685 27.300 65.945 27.800 ;
        RECT 68.965 27.300 69.225 27.800 ;
        RECT 72.245 27.300 72.505 27.800 ;
        RECT 79.525 27.300 79.785 27.800 ;
        RECT 86.805 27.300 87.065 27.800 ;
        RECT 90.085 27.300 90.345 27.800 ;
        RECT 93.365 27.300 93.625 27.800 ;
        RECT 94.380 27.110 94.670 27.990 ;
        RECT 64.640 26.820 72.115 27.110 ;
        RECT 87.205 26.820 94.670 27.110 ;
        RECT 64.640 25.540 64.930 26.820 ;
        RECT 94.380 25.540 94.670 26.820 ;
        RECT 124.750 26.555 125.040 29.625 ;
        RECT 125.700 29.585 126.290 29.625 ;
        RECT 126.560 29.585 128.010 29.915 ;
        RECT 128.280 29.625 129.820 29.915 ;
        RECT 128.280 29.585 128.870 29.625 ;
        RECT 125.450 29.245 125.680 29.395 ;
        RECT 125.880 29.245 126.110 29.395 ;
        RECT 126.310 29.245 126.540 29.395 ;
        RECT 125.435 28.395 125.695 29.245 ;
        RECT 125.865 28.395 126.125 29.245 ;
        RECT 126.295 28.395 126.555 29.245 ;
        RECT 126.725 28.395 126.985 29.395 ;
        RECT 127.170 29.245 127.400 29.395 ;
        RECT 127.155 28.395 127.415 29.245 ;
        RECT 127.585 28.395 127.845 29.395 ;
        RECT 128.030 29.245 128.260 29.395 ;
        RECT 128.460 29.245 128.690 29.395 ;
        RECT 128.890 29.245 129.120 29.395 ;
        RECT 129.530 29.245 129.820 29.625 ;
        RECT 128.015 28.395 128.275 29.245 ;
        RECT 128.445 28.395 128.705 29.245 ;
        RECT 128.875 28.395 129.135 29.245 ;
        RECT 129.525 28.395 129.820 29.245 ;
        RECT 125.450 27.670 125.680 27.745 ;
        RECT 125.880 27.670 126.110 27.745 ;
        RECT 125.435 26.820 125.695 27.670 ;
        RECT 125.865 26.820 126.125 27.670 ;
        RECT 125.450 26.745 125.680 26.820 ;
        RECT 125.880 26.745 126.110 26.820 ;
        RECT 126.295 26.745 126.555 27.745 ;
        RECT 126.725 26.745 126.985 27.745 ;
        RECT 127.155 26.745 127.415 27.745 ;
        RECT 127.585 26.745 127.845 27.745 ;
        RECT 128.015 26.745 128.275 27.745 ;
        RECT 128.460 27.670 128.690 27.745 ;
        RECT 128.890 27.670 129.120 27.745 ;
        RECT 129.530 27.670 129.820 28.395 ;
        RECT 135.060 34.270 135.350 34.820 ;
        RECT 135.755 34.800 137.745 35.130 ;
        RECT 137.415 34.270 137.745 34.800 ;
        RECT 137.885 35.130 138.165 35.445 ;
        RECT 140.440 35.130 140.770 35.660 ;
        RECT 137.885 34.800 140.770 35.130 ;
        RECT 144.140 35.110 144.430 35.660 ;
        RECT 137.885 34.485 138.165 34.800 ;
        RECT 140.440 34.270 140.770 34.800 ;
        RECT 144.140 34.270 144.430 34.820 ;
        RECT 135.060 33.980 136.600 34.270 ;
        RECT 136.870 33.980 138.320 34.270 ;
        RECT 138.590 33.980 142.620 34.270 ;
        RECT 142.890 33.980 144.430 34.270 ;
        RECT 135.060 31.390 135.350 33.980 ;
        RECT 135.760 33.290 135.990 33.790 ;
        RECT 136.190 33.290 136.420 33.790 ;
        RECT 136.620 33.290 136.850 33.790 ;
        RECT 135.745 32.290 136.005 33.290 ;
        RECT 136.175 32.290 136.435 33.290 ;
        RECT 136.605 32.290 136.865 33.290 ;
        RECT 135.760 31.790 135.990 32.290 ;
        RECT 136.190 31.790 136.420 32.290 ;
        RECT 136.620 31.790 136.850 32.290 ;
        RECT 137.035 31.790 137.295 33.790 ;
        RECT 137.480 33.290 137.710 33.790 ;
        RECT 137.465 32.290 137.725 33.290 ;
        RECT 137.480 31.790 137.710 32.290 ;
        RECT 137.895 31.790 138.155 33.790 ;
        RECT 138.340 33.290 138.570 33.790 ;
        RECT 138.325 32.290 138.585 33.290 ;
        RECT 138.340 31.790 138.570 32.290 ;
        RECT 138.755 31.790 139.015 33.790 ;
        RECT 139.200 33.290 139.430 33.790 ;
        RECT 139.185 32.290 139.445 33.290 ;
        RECT 139.200 31.790 139.430 32.290 ;
        RECT 139.615 31.790 139.875 33.790 ;
        RECT 140.060 33.290 140.290 33.790 ;
        RECT 140.045 32.290 140.305 33.290 ;
        RECT 140.060 31.790 140.290 32.290 ;
        RECT 140.475 31.790 140.735 33.790 ;
        RECT 140.920 33.290 141.150 33.790 ;
        RECT 140.905 32.290 141.165 33.290 ;
        RECT 140.920 31.790 141.150 32.290 ;
        RECT 141.335 31.790 141.595 33.790 ;
        RECT 141.780 33.290 142.010 33.790 ;
        RECT 141.765 32.290 142.025 33.290 ;
        RECT 141.780 31.790 142.010 32.290 ;
        RECT 142.195 31.790 142.455 33.790 ;
        RECT 142.640 33.290 142.870 33.790 ;
        RECT 143.070 33.290 143.300 33.790 ;
        RECT 143.500 33.290 143.730 33.790 ;
        RECT 142.625 32.290 142.885 33.290 ;
        RECT 143.055 32.290 143.315 33.290 ;
        RECT 143.485 32.290 143.745 33.290 ;
        RECT 142.640 31.790 142.870 32.290 ;
        RECT 143.070 31.790 143.300 32.290 ;
        RECT 143.500 31.790 143.730 32.290 ;
        RECT 144.140 31.390 144.430 33.980 ;
        RECT 135.060 31.100 144.430 31.390 ;
        RECT 135.060 28.510 135.350 31.100 ;
        RECT 135.760 30.200 135.990 30.700 ;
        RECT 136.190 30.200 136.420 30.700 ;
        RECT 136.620 30.200 136.850 30.700 ;
        RECT 135.745 29.200 136.005 30.200 ;
        RECT 136.175 29.200 136.435 30.200 ;
        RECT 136.605 29.200 136.865 30.200 ;
        RECT 135.760 28.700 135.990 29.200 ;
        RECT 136.190 28.700 136.420 29.200 ;
        RECT 136.620 28.700 136.850 29.200 ;
        RECT 137.035 28.700 137.295 30.700 ;
        RECT 137.480 30.200 137.710 30.700 ;
        RECT 137.465 29.200 137.725 30.200 ;
        RECT 137.480 28.700 137.710 29.200 ;
        RECT 137.895 28.700 138.155 30.700 ;
        RECT 138.340 30.200 138.570 30.700 ;
        RECT 138.325 29.200 138.585 30.200 ;
        RECT 138.340 28.700 138.570 29.200 ;
        RECT 138.755 28.700 139.015 30.700 ;
        RECT 139.200 30.200 139.430 30.700 ;
        RECT 139.185 29.200 139.445 30.200 ;
        RECT 139.200 28.700 139.430 29.200 ;
        RECT 139.615 28.700 139.875 30.700 ;
        RECT 140.060 30.200 140.290 30.700 ;
        RECT 140.045 29.200 140.305 30.200 ;
        RECT 140.060 28.700 140.290 29.200 ;
        RECT 140.475 28.700 140.735 30.700 ;
        RECT 140.920 30.200 141.150 30.700 ;
        RECT 140.905 29.200 141.165 30.200 ;
        RECT 140.920 28.700 141.150 29.200 ;
        RECT 141.335 28.700 141.595 30.700 ;
        RECT 141.780 30.200 142.010 30.700 ;
        RECT 141.765 29.200 142.025 30.200 ;
        RECT 141.780 28.700 142.010 29.200 ;
        RECT 142.195 28.700 142.455 30.700 ;
        RECT 142.640 30.200 142.870 30.700 ;
        RECT 143.070 30.200 143.300 30.700 ;
        RECT 143.500 30.200 143.730 30.700 ;
        RECT 142.625 29.200 142.885 30.200 ;
        RECT 143.055 29.200 143.315 30.200 ;
        RECT 143.485 29.200 143.745 30.200 ;
        RECT 142.640 28.700 142.870 29.200 ;
        RECT 143.070 28.700 143.300 29.200 ;
        RECT 143.500 28.700 143.730 29.200 ;
        RECT 144.140 28.510 144.430 31.100 ;
        RECT 135.060 28.220 136.600 28.510 ;
        RECT 136.870 28.220 138.320 28.510 ;
        RECT 138.590 28.220 142.620 28.510 ;
        RECT 142.890 28.220 144.430 28.510 ;
        RECT 135.060 27.670 135.350 28.220 ;
        RECT 137.415 27.690 137.745 28.220 ;
        RECT 128.445 26.820 128.705 27.670 ;
        RECT 128.875 26.820 129.135 27.670 ;
        RECT 129.525 26.820 129.820 27.670 ;
        RECT 128.460 26.745 128.690 26.820 ;
        RECT 128.890 26.745 129.120 26.820 ;
        RECT 129.530 26.555 129.820 26.820 ;
        RECT 124.750 26.265 126.290 26.555 ;
        RECT 124.750 25.800 125.040 26.265 ;
        RECT 126.560 26.225 128.010 26.555 ;
        RECT 128.280 26.265 129.820 26.555 ;
        RECT 127.550 25.760 127.880 26.225 ;
        RECT 129.530 25.800 129.820 26.265 ;
        RECT 135.060 26.830 135.350 27.380 ;
        RECT 135.755 27.360 137.745 27.690 ;
        RECT 137.415 26.830 137.745 27.360 ;
        RECT 137.885 27.690 138.165 28.005 ;
        RECT 140.440 27.690 140.770 28.220 ;
        RECT 137.885 27.360 140.770 27.690 ;
        RECT 144.140 27.670 144.430 28.220 ;
        RECT 137.885 27.045 138.165 27.360 ;
        RECT 140.440 26.830 140.770 27.360 ;
        RECT 144.140 26.830 144.430 27.380 ;
        RECT 135.060 26.540 136.600 26.830 ;
        RECT 136.870 26.540 138.320 26.830 ;
        RECT 138.590 26.540 142.620 26.830 ;
        RECT 142.890 26.540 144.430 26.830 ;
        RECT 64.640 25.250 67.715 25.540 ;
        RECT 68.280 25.250 69.950 25.540 ;
        RECT 70.560 25.250 72.230 25.540 ;
        RECT 72.840 25.250 74.510 25.540 ;
        RECT 75.120 25.250 76.790 25.540 ;
        RECT 77.365 25.250 81.955 25.540 ;
        RECT 82.520 25.250 84.190 25.540 ;
        RECT 84.800 25.250 86.470 25.540 ;
        RECT 87.080 25.250 88.750 25.540 ;
        RECT 89.360 25.250 91.030 25.540 ;
        RECT 91.605 25.250 94.670 25.540 ;
        RECT 125.505 25.430 127.880 25.760 ;
        RECT 64.640 23.820 64.930 25.250 ;
        RECT 65.285 24.560 65.545 25.060 ;
        RECT 66.580 24.560 66.810 25.250 ;
        RECT 67.845 24.560 68.105 25.060 ;
        RECT 70.125 24.560 70.385 25.060 ;
        RECT 72.405 24.560 72.665 25.060 ;
        RECT 74.685 24.560 74.945 25.060 ;
        RECT 76.965 24.560 77.225 25.060 ;
        RECT 78.235 24.370 78.515 25.250 ;
        RECT 79.515 24.370 79.795 25.250 ;
        RECT 80.795 24.370 81.075 25.250 ;
        RECT 82.085 24.560 82.345 25.060 ;
        RECT 84.365 24.560 84.625 25.060 ;
        RECT 86.645 24.560 86.905 25.060 ;
        RECT 88.925 24.560 89.185 25.060 ;
        RECT 91.205 24.560 91.465 25.060 ;
        RECT 92.500 24.560 92.730 25.250 ;
        RECT 93.765 24.560 94.025 25.060 ;
        RECT 66.280 24.040 76.790 24.370 ;
        RECT 77.365 24.080 81.955 24.370 ;
        RECT 82.520 24.040 93.030 24.370 ;
        RECT 94.380 23.820 94.670 25.250 ;
        RECT 64.640 23.530 94.670 23.820 ;
        RECT 124.750 24.925 125.040 25.390 ;
        RECT 127.550 24.925 127.880 25.430 ;
        RECT 129.530 24.925 129.820 25.390 ;
        RECT 124.750 24.635 126.290 24.925 ;
        RECT 126.560 24.635 127.150 24.925 ;
        RECT 127.420 24.635 128.010 24.925 ;
        RECT 128.280 24.635 129.820 24.925 ;
        RECT 135.060 24.975 135.350 26.540 ;
        RECT 135.745 25.350 136.005 26.350 ;
        RECT 136.175 25.350 136.435 26.350 ;
        RECT 136.605 25.350 136.865 26.350 ;
        RECT 137.035 25.350 137.295 26.350 ;
        RECT 137.465 25.350 137.725 26.350 ;
        RECT 137.895 25.350 138.155 26.350 ;
        RECT 138.325 25.350 138.585 26.350 ;
        RECT 138.755 25.350 139.015 26.350 ;
        RECT 139.185 25.350 139.445 26.350 ;
        RECT 139.615 25.350 139.875 26.350 ;
        RECT 140.045 25.350 140.305 26.350 ;
        RECT 140.475 25.350 140.735 26.350 ;
        RECT 140.905 25.350 141.165 26.350 ;
        RECT 141.335 25.350 141.595 26.350 ;
        RECT 141.765 25.350 142.025 26.350 ;
        RECT 142.195 25.350 142.455 26.350 ;
        RECT 142.625 25.350 142.885 26.350 ;
        RECT 143.055 25.350 143.315 26.350 ;
        RECT 143.485 25.350 143.745 26.350 ;
        RECT 144.140 24.975 144.430 26.540 ;
        RECT 135.060 24.685 144.430 24.975 ;
        RECT 124.750 22.705 125.040 24.635 ;
        RECT 129.530 24.445 129.820 24.635 ;
        RECT 125.435 23.595 125.695 24.445 ;
        RECT 125.865 23.595 126.125 24.445 ;
        RECT 126.295 23.595 126.555 24.445 ;
        RECT 125.450 23.445 125.680 23.595 ;
        RECT 125.880 23.445 126.110 23.595 ;
        RECT 126.310 23.445 126.540 23.595 ;
        RECT 126.725 23.445 126.985 24.445 ;
        RECT 127.155 23.595 127.415 24.445 ;
        RECT 127.170 23.445 127.400 23.595 ;
        RECT 127.585 23.445 127.845 24.445 ;
        RECT 128.015 23.595 128.275 24.445 ;
        RECT 128.445 23.595 128.705 24.445 ;
        RECT 128.875 23.595 129.135 24.445 ;
        RECT 129.525 23.595 129.820 24.445 ;
        RECT 128.030 23.445 128.260 23.595 ;
        RECT 128.460 23.445 128.690 23.595 ;
        RECT 128.890 23.445 129.120 23.595 ;
        RECT 125.700 22.965 126.290 23.255 ;
        RECT 126.560 22.925 127.150 23.255 ;
        RECT 127.420 22.965 128.010 23.255 ;
        RECT 128.280 22.965 128.870 23.255 ;
        RECT 129.530 22.705 129.820 23.595 ;
        RECT 124.750 22.415 129.820 22.705 ;
        RECT 69.130 21.900 90.120 22.190 ;
        RECT 69.130 21.620 69.420 21.900 ;
        RECT 70.215 21.620 72.245 21.640 ;
        RECT 69.130 21.330 72.245 21.620 ;
        RECT 72.810 21.330 76.760 21.660 ;
        RECT 77.335 21.620 79.365 21.640 ;
        RECT 79.895 21.620 81.925 21.640 ;
        RECT 77.335 21.330 81.925 21.620 ;
        RECT 82.490 21.330 86.440 21.660 ;
        RECT 87.015 21.620 89.045 21.640 ;
        RECT 89.830 21.620 90.120 21.900 ;
        RECT 87.015 21.330 90.120 21.620 ;
        RECT 69.130 19.990 69.420 21.330 ;
        RECT 69.815 20.160 70.075 21.160 ;
        RECT 71.095 20.160 71.355 21.160 ;
        RECT 72.375 20.160 72.635 21.160 ;
        RECT 74.670 20.160 74.935 21.330 ;
        RECT 76.935 20.160 77.195 21.160 ;
        RECT 78.205 19.990 78.485 21.330 ;
        RECT 79.485 19.990 79.765 21.330 ;
        RECT 80.765 19.990 81.045 21.330 ;
        RECT 82.055 20.160 82.315 21.160 ;
        RECT 84.350 20.160 84.625 21.330 ;
        RECT 86.615 20.160 86.875 21.160 ;
        RECT 87.895 20.160 88.155 21.160 ;
        RECT 89.175 20.160 89.435 21.160 ;
        RECT 89.830 19.990 90.120 21.330 ;
        RECT 135.060 22.080 144.430 22.370 ;
        RECT 69.130 19.700 72.245 19.990 ;
        RECT 69.130 19.420 69.420 19.700 ;
        RECT 70.215 19.680 72.245 19.700 ;
        RECT 72.810 19.640 76.760 19.970 ;
        RECT 77.335 19.700 81.925 19.990 ;
        RECT 77.335 19.680 79.365 19.700 ;
        RECT 79.895 19.680 81.925 19.700 ;
        RECT 87.015 19.700 90.120 19.990 ;
        RECT 87.015 19.680 89.045 19.700 ;
        RECT 89.830 19.420 90.120 19.700 ;
        RECT 69.130 19.130 90.120 19.420 ;
        RECT 94.080 21.015 118.510 21.305 ;
        RECT 94.080 19.925 94.370 21.015 ;
        RECT 94.765 20.115 95.025 20.615 ;
        RECT 97.045 20.115 97.305 20.615 ;
        RECT 99.325 20.115 99.585 20.615 ;
        RECT 101.605 20.115 101.865 20.615 ;
        RECT 103.885 20.115 104.145 20.615 ;
        RECT 106.165 20.115 106.425 20.615 ;
        RECT 108.445 20.115 108.705 20.615 ;
        RECT 110.725 20.115 110.985 20.615 ;
        RECT 113.005 20.115 113.265 20.615 ;
        RECT 115.285 20.115 115.545 20.615 ;
        RECT 117.565 20.115 117.825 20.615 ;
        RECT 118.220 19.925 118.510 21.015 ;
        RECT 94.080 19.635 99.150 19.925 ;
        RECT 94.080 18.610 94.370 19.635 ;
        RECT 99.760 19.595 103.710 19.925 ;
        RECT 104.320 19.595 108.270 19.925 ;
        RECT 108.880 19.595 112.830 19.925 ;
        RECT 113.440 19.635 118.510 19.925 ;
        RECT 101.595 18.670 101.875 18.985 ;
        RECT 104.320 18.670 104.650 19.595 ;
        RECT 55.920 17.645 65.230 17.935 ;
        RECT 55.920 17.385 56.210 17.645 ;
        RECT 64.940 17.385 65.230 17.645 ;
        RECT 55.920 17.095 57.990 17.385 ;
        RECT 63.160 17.095 65.230 17.385 ;
        RECT 55.920 15.665 56.210 17.095 ;
        RECT 56.605 16.405 56.865 16.905 ;
        RECT 57.385 16.405 57.645 16.905 ;
        RECT 58.165 16.405 58.425 16.905 ;
        RECT 60.445 16.405 60.705 16.905 ;
        RECT 62.725 16.405 62.985 16.905 ;
        RECT 63.505 16.405 63.765 16.905 ;
        RECT 64.285 16.405 64.545 16.905 ;
        RECT 58.600 15.885 62.550 16.215 ;
        RECT 64.940 15.665 65.230 17.095 ;
        RECT 55.920 15.375 65.230 15.665 ;
        RECT 69.130 17.645 90.120 17.935 ;
        RECT 69.130 17.365 69.420 17.645 ;
        RECT 70.215 17.365 72.245 17.385 ;
        RECT 69.130 17.075 72.245 17.365 ;
        RECT 72.810 17.095 76.760 17.425 ;
        RECT 77.335 17.365 79.365 17.385 ;
        RECT 79.895 17.365 81.925 17.385 ;
        RECT 69.130 16.215 69.420 17.075 ;
        RECT 69.815 16.405 70.075 16.905 ;
        RECT 71.095 16.405 71.355 16.905 ;
        RECT 72.375 16.405 72.635 16.905 ;
        RECT 74.635 16.215 74.925 17.095 ;
        RECT 77.335 17.075 81.925 17.365 ;
        RECT 87.015 17.365 89.045 17.385 ;
        RECT 89.830 17.365 90.120 17.645 ;
        RECT 87.015 17.075 90.120 17.365 ;
        RECT 76.935 16.405 77.195 16.905 ;
        RECT 78.205 16.215 78.485 17.075 ;
        RECT 79.485 16.215 79.765 17.075 ;
        RECT 80.765 16.215 81.045 17.075 ;
        RECT 82.055 16.405 82.315 16.905 ;
        RECT 84.335 16.405 84.595 16.905 ;
        RECT 86.615 16.405 86.875 16.905 ;
        RECT 87.895 16.405 88.155 16.905 ;
        RECT 89.175 16.405 89.435 16.905 ;
        RECT 89.830 16.215 90.120 17.075 ;
        RECT 69.130 15.925 72.245 16.215 ;
        RECT 69.130 15.665 69.420 15.925 ;
        RECT 72.675 15.885 76.760 16.215 ;
        RECT 77.335 15.925 81.925 16.215 ;
        RECT 82.490 16.210 84.160 16.215 ;
        RECT 84.770 16.210 86.440 16.215 ;
        RECT 82.490 15.880 86.440 16.210 ;
        RECT 87.015 15.925 90.120 16.215 ;
        RECT 89.830 15.665 90.120 15.925 ;
        RECT 69.130 15.375 90.120 15.665 ;
        RECT 94.080 16.795 94.370 18.345 ;
        RECT 101.595 18.340 104.650 18.670 ;
        RECT 101.595 18.025 101.875 18.340 ;
        RECT 104.320 16.835 104.650 18.340 ;
        RECT 106.155 18.670 106.435 18.985 ;
        RECT 108.880 18.670 109.210 19.595 ;
        RECT 106.155 18.340 109.210 18.670 ;
        RECT 118.220 18.610 118.510 19.635 ;
        RECT 135.060 19.490 135.350 22.080 ;
        RECT 135.760 21.180 135.990 21.680 ;
        RECT 136.190 21.180 136.420 21.680 ;
        RECT 136.620 21.180 136.850 21.680 ;
        RECT 135.745 20.180 136.005 21.180 ;
        RECT 136.175 20.180 136.435 21.180 ;
        RECT 136.605 20.180 136.865 21.180 ;
        RECT 135.760 19.680 135.990 20.180 ;
        RECT 136.190 19.680 136.420 20.180 ;
        RECT 136.620 19.680 136.850 20.180 ;
        RECT 137.035 19.680 137.295 21.680 ;
        RECT 137.480 21.180 137.710 21.680 ;
        RECT 137.465 20.180 137.725 21.180 ;
        RECT 137.480 19.680 137.710 20.180 ;
        RECT 137.895 19.680 138.155 21.680 ;
        RECT 138.340 21.180 138.570 21.680 ;
        RECT 138.325 20.180 138.585 21.180 ;
        RECT 138.340 19.680 138.570 20.180 ;
        RECT 138.755 19.680 139.015 21.680 ;
        RECT 139.200 21.180 139.430 21.680 ;
        RECT 139.185 20.180 139.445 21.180 ;
        RECT 139.200 19.680 139.430 20.180 ;
        RECT 139.615 19.680 139.875 21.680 ;
        RECT 140.060 21.180 140.290 21.680 ;
        RECT 140.045 20.180 140.305 21.180 ;
        RECT 140.060 19.680 140.290 20.180 ;
        RECT 140.475 19.680 140.735 21.680 ;
        RECT 140.920 21.180 141.150 21.680 ;
        RECT 140.905 20.180 141.165 21.180 ;
        RECT 140.920 19.680 141.150 20.180 ;
        RECT 141.335 19.680 141.595 21.680 ;
        RECT 141.780 21.180 142.010 21.680 ;
        RECT 141.765 20.180 142.025 21.180 ;
        RECT 141.780 19.680 142.010 20.180 ;
        RECT 142.195 19.680 142.455 21.680 ;
        RECT 142.640 21.180 142.870 21.680 ;
        RECT 143.070 21.180 143.300 21.680 ;
        RECT 143.500 21.180 143.730 21.680 ;
        RECT 142.625 20.180 142.885 21.180 ;
        RECT 143.055 20.180 143.315 21.180 ;
        RECT 143.485 20.180 143.745 21.180 ;
        RECT 142.640 19.680 142.870 20.180 ;
        RECT 143.070 19.680 143.300 20.180 ;
        RECT 143.500 19.680 143.730 20.180 ;
        RECT 144.140 19.490 144.430 22.080 ;
        RECT 135.060 19.200 136.600 19.490 ;
        RECT 136.870 19.200 138.320 19.490 ;
        RECT 138.590 19.200 142.620 19.490 ;
        RECT 142.890 19.200 144.430 19.490 ;
        RECT 135.060 18.650 135.350 19.200 ;
        RECT 137.415 18.670 137.745 19.200 ;
        RECT 106.155 18.025 106.435 18.340 ;
        RECT 108.880 16.835 109.210 18.340 ;
        RECT 94.080 16.505 99.150 16.795 ;
        RECT 99.760 16.505 103.710 16.835 ;
        RECT 104.320 16.505 108.270 16.835 ;
        RECT 108.880 16.505 112.830 16.835 ;
        RECT 118.220 16.795 118.510 18.345 ;
        RECT 113.440 16.505 118.510 16.795 ;
        RECT 94.080 14.915 94.370 16.505 ;
        RECT 94.765 15.315 95.025 16.315 ;
        RECT 97.045 15.315 97.305 16.315 ;
        RECT 99.325 15.315 99.585 16.315 ;
        RECT 101.605 15.315 101.865 16.315 ;
        RECT 103.885 15.315 104.145 16.315 ;
        RECT 106.165 15.315 106.425 16.315 ;
        RECT 108.445 15.315 108.705 16.315 ;
        RECT 110.725 15.315 110.985 16.315 ;
        RECT 113.005 15.315 113.265 16.315 ;
        RECT 115.285 15.315 115.545 16.315 ;
        RECT 117.565 15.315 117.825 16.315 ;
        RECT 118.220 14.915 118.510 16.505 ;
        RECT 135.060 17.810 135.350 18.360 ;
        RECT 135.755 18.340 137.745 18.670 ;
        RECT 137.415 17.810 137.745 18.340 ;
        RECT 137.885 18.670 138.165 18.985 ;
        RECT 140.440 18.670 140.770 19.200 ;
        RECT 137.885 18.340 140.770 18.670 ;
        RECT 144.140 18.650 144.430 19.200 ;
        RECT 137.885 18.025 138.165 18.340 ;
        RECT 140.440 17.810 140.770 18.340 ;
        RECT 144.140 17.810 144.430 18.360 ;
        RECT 135.060 17.520 136.600 17.810 ;
        RECT 136.870 17.520 138.320 17.810 ;
        RECT 138.590 17.520 142.620 17.810 ;
        RECT 142.890 17.520 144.430 17.810 ;
        RECT 135.060 15.955 135.350 17.520 ;
        RECT 135.745 16.330 136.005 17.330 ;
        RECT 136.175 16.330 136.435 17.330 ;
        RECT 136.605 16.330 136.865 17.330 ;
        RECT 137.035 16.330 137.295 17.330 ;
        RECT 137.465 16.330 137.725 17.330 ;
        RECT 137.895 16.330 138.155 17.330 ;
        RECT 138.325 16.330 138.585 17.330 ;
        RECT 138.755 16.330 139.015 17.330 ;
        RECT 139.185 16.330 139.445 17.330 ;
        RECT 139.615 16.330 139.875 17.330 ;
        RECT 140.045 16.330 140.305 17.330 ;
        RECT 140.475 16.330 140.735 17.330 ;
        RECT 140.905 16.330 141.165 17.330 ;
        RECT 141.335 16.330 141.595 17.330 ;
        RECT 141.765 16.330 142.025 17.330 ;
        RECT 142.195 16.330 142.455 17.330 ;
        RECT 142.625 16.330 142.885 17.330 ;
        RECT 143.055 16.330 143.315 17.330 ;
        RECT 143.485 16.330 143.745 17.330 ;
        RECT 144.140 15.955 144.430 17.520 ;
        RECT 135.060 15.665 144.430 15.955 ;
        RECT 94.080 14.625 118.510 14.915 ;
        RECT 55.920 13.480 95.710 13.770 ;
        RECT 55.920 11.550 56.210 13.480 ;
        RECT 58.600 12.930 62.550 13.260 ;
        RECT 66.280 12.930 79.350 13.260 ;
        RECT 79.960 12.930 93.030 13.260 ;
        RECT 56.605 11.740 56.865 12.740 ;
        RECT 57.385 11.740 57.645 12.740 ;
        RECT 58.165 11.740 58.425 12.740 ;
        RECT 60.445 11.740 60.705 12.740 ;
        RECT 62.725 11.740 62.985 12.740 ;
        RECT 63.490 11.550 63.780 12.740 ;
        RECT 64.270 11.550 64.560 12.740 ;
        RECT 65.050 11.550 65.340 12.740 ;
        RECT 65.845 11.740 66.105 12.740 ;
        RECT 68.125 11.740 68.385 12.740 ;
        RECT 70.405 11.740 70.665 12.740 ;
        RECT 72.685 11.740 72.945 12.740 ;
        RECT 74.965 11.740 75.225 12.740 ;
        RECT 77.245 11.740 77.505 12.740 ;
        RECT 79.525 11.740 79.785 12.740 ;
        RECT 81.805 11.740 82.065 12.740 ;
        RECT 84.085 11.740 84.345 12.740 ;
        RECT 86.365 11.740 86.625 12.740 ;
        RECT 88.645 11.740 88.905 12.740 ;
        RECT 90.925 11.740 91.185 12.740 ;
        RECT 93.205 11.740 93.465 12.740 ;
        RECT 93.985 11.740 94.245 12.740 ;
        RECT 94.765 11.740 95.025 12.740 ;
        RECT 95.420 11.550 95.710 13.480 ;
        RECT 55.920 11.260 57.990 11.550 ;
        RECT 63.160 11.260 65.670 11.550 ;
        RECT 66.280 11.260 67.950 11.550 ;
        RECT 68.560 11.260 70.230 11.550 ;
        RECT 70.840 11.260 72.510 11.550 ;
        RECT 73.120 11.260 74.790 11.550 ;
        RECT 75.400 11.260 77.070 11.550 ;
        RECT 77.680 11.260 79.350 11.550 ;
        RECT 79.960 11.260 81.630 11.550 ;
        RECT 82.240 11.260 83.910 11.550 ;
        RECT 84.520 11.260 86.190 11.550 ;
        RECT 86.800 11.260 88.470 11.550 ;
        RECT 89.080 11.260 90.750 11.550 ;
        RECT 91.360 11.260 93.030 11.550 ;
        RECT 93.640 11.260 95.710 11.550 ;
        RECT 55.920 9.630 56.210 11.260 ;
        RECT 95.420 9.630 95.710 11.260 ;
        RECT 55.920 9.340 77.070 9.630 ;
        RECT 82.240 9.340 95.710 9.630 ;
        RECT 55.920 7.410 56.210 9.340 ;
        RECT 65.845 8.150 66.105 9.150 ;
        RECT 68.125 8.150 68.385 9.150 ;
        RECT 70.405 8.150 70.665 9.150 ;
        RECT 72.685 8.150 72.945 9.150 ;
        RECT 74.965 8.150 75.225 9.150 ;
        RECT 77.245 8.150 77.505 9.150 ;
        RECT 79.525 8.150 79.785 9.150 ;
        RECT 81.805 8.150 82.065 9.150 ;
        RECT 84.085 8.150 84.345 9.150 ;
        RECT 86.365 8.150 86.625 9.150 ;
        RECT 88.645 8.150 88.905 9.150 ;
        RECT 90.925 8.150 91.185 9.150 ;
        RECT 93.205 8.150 93.465 9.150 ;
        RECT 77.680 7.630 81.630 7.960 ;
        RECT 95.420 7.410 95.710 9.340 ;
        RECT 55.920 7.120 95.710 7.410 ;
      LAYER via ;
        RECT 141.750 77.335 142.010 77.595 ;
        RECT 142.070 77.335 142.330 77.595 ;
        RECT 142.390 77.335 142.650 77.595 ;
        RECT 42.725 75.560 42.985 75.820 ;
        RECT 42.725 75.240 42.985 75.500 ;
        RECT 43.355 75.560 43.615 75.820 ;
        RECT 43.355 75.240 43.615 75.500 ;
        RECT 45.635 75.560 45.895 75.820 ;
        RECT 45.635 75.240 45.895 75.500 ;
        RECT 47.915 75.560 48.175 75.820 ;
        RECT 47.915 75.240 48.175 75.500 ;
        RECT 50.195 75.560 50.455 75.820 ;
        RECT 50.195 75.240 50.455 75.500 ;
        RECT 52.475 75.560 52.735 75.820 ;
        RECT 52.475 75.240 52.735 75.500 ;
        RECT 54.755 75.560 55.015 75.820 ;
        RECT 54.755 75.240 55.015 75.500 ;
        RECT 57.035 75.560 57.295 75.820 ;
        RECT 57.035 75.240 57.295 75.500 ;
        RECT 59.315 75.560 59.575 75.820 ;
        RECT 59.315 75.240 59.575 75.500 ;
        RECT 61.595 75.560 61.855 75.820 ;
        RECT 61.595 75.240 61.855 75.500 ;
        RECT 63.875 75.560 64.135 75.820 ;
        RECT 63.875 75.240 64.135 75.500 ;
        RECT 66.155 75.560 66.415 75.820 ;
        RECT 66.155 75.240 66.415 75.500 ;
        RECT 68.435 75.560 68.695 75.820 ;
        RECT 68.435 75.240 68.695 75.500 ;
        RECT 70.715 75.560 70.975 75.820 ;
        RECT 70.715 75.240 70.975 75.500 ;
        RECT 72.995 75.560 73.255 75.820 ;
        RECT 72.995 75.240 73.255 75.500 ;
        RECT 75.275 75.560 75.535 75.820 ;
        RECT 75.275 75.240 75.535 75.500 ;
        RECT 77.555 75.560 77.815 75.820 ;
        RECT 77.555 75.240 77.815 75.500 ;
        RECT 79.835 75.560 80.095 75.820 ;
        RECT 79.835 75.240 80.095 75.500 ;
        RECT 82.115 75.560 82.375 75.820 ;
        RECT 82.115 75.240 82.375 75.500 ;
        RECT 84.395 75.560 84.655 75.820 ;
        RECT 84.395 75.240 84.655 75.500 ;
        RECT 86.675 75.560 86.935 75.820 ;
        RECT 86.675 75.240 86.935 75.500 ;
        RECT 88.955 75.560 89.215 75.820 ;
        RECT 88.955 75.240 89.215 75.500 ;
        RECT 91.235 75.560 91.495 75.820 ;
        RECT 91.235 75.240 91.495 75.500 ;
        RECT 93.515 75.560 93.775 75.820 ;
        RECT 93.515 75.240 93.775 75.500 ;
        RECT 95.795 75.560 96.055 75.820 ;
        RECT 95.795 75.240 96.055 75.500 ;
        RECT 98.075 75.560 98.335 75.820 ;
        RECT 98.075 75.240 98.335 75.500 ;
        RECT 100.355 75.560 100.615 75.820 ;
        RECT 100.355 75.240 100.615 75.500 ;
        RECT 102.635 75.560 102.895 75.820 ;
        RECT 102.635 75.240 102.895 75.500 ;
        RECT 104.915 75.560 105.175 75.820 ;
        RECT 104.915 75.240 105.175 75.500 ;
        RECT 107.195 75.560 107.455 75.820 ;
        RECT 107.195 75.240 107.455 75.500 ;
        RECT 109.475 75.560 109.735 75.820 ;
        RECT 109.475 75.240 109.735 75.500 ;
        RECT 111.755 75.560 112.015 75.820 ;
        RECT 111.755 75.240 112.015 75.500 ;
        RECT 114.035 75.560 114.295 75.820 ;
        RECT 114.035 75.240 114.295 75.500 ;
        RECT 116.315 75.560 116.575 75.820 ;
        RECT 116.315 75.240 116.575 75.500 ;
        RECT 118.595 75.560 118.855 75.820 ;
        RECT 118.595 75.240 118.855 75.500 ;
        RECT 120.875 75.560 121.135 75.820 ;
        RECT 120.875 75.240 121.135 75.500 ;
        RECT 123.155 75.560 123.415 75.820 ;
        RECT 123.155 75.240 123.415 75.500 ;
        RECT 125.435 75.560 125.695 75.820 ;
        RECT 125.435 75.240 125.695 75.500 ;
        RECT 127.715 75.560 127.975 75.820 ;
        RECT 127.715 75.240 127.975 75.500 ;
        RECT 129.995 75.560 130.255 75.820 ;
        RECT 129.995 75.240 130.255 75.500 ;
        RECT 130.625 75.560 130.885 75.820 ;
        RECT 130.625 75.240 130.885 75.500 ;
        RECT 137.125 76.805 137.385 77.065 ;
        RECT 137.125 76.485 137.385 76.745 ;
        RECT 137.755 76.805 138.015 77.065 ;
        RECT 137.755 76.485 138.015 76.745 ;
        RECT 138.185 76.805 138.445 77.065 ;
        RECT 138.185 76.485 138.445 76.745 ;
        RECT 138.615 76.805 138.875 77.065 ;
        RECT 138.615 76.485 138.875 76.745 ;
        RECT 139.045 76.805 139.305 77.065 ;
        RECT 139.045 76.485 139.305 76.745 ;
        RECT 139.475 76.805 139.735 77.065 ;
        RECT 139.475 76.485 139.735 76.745 ;
        RECT 139.905 76.805 140.165 77.065 ;
        RECT 139.905 76.485 140.165 76.745 ;
        RECT 140.335 76.805 140.595 77.065 ;
        RECT 140.335 76.485 140.595 76.745 ;
        RECT 140.765 76.805 141.025 77.065 ;
        RECT 140.765 76.485 141.025 76.745 ;
        RECT 141.195 76.805 141.455 77.065 ;
        RECT 141.195 76.485 141.455 76.745 ;
        RECT 141.625 76.805 141.885 77.065 ;
        RECT 141.625 76.485 141.885 76.745 ;
        RECT 142.055 76.805 142.315 77.065 ;
        RECT 142.055 76.485 142.315 76.745 ;
        RECT 142.485 76.805 142.745 77.065 ;
        RECT 142.485 76.485 142.745 76.745 ;
        RECT 142.915 76.805 143.175 77.065 ;
        RECT 142.915 76.485 143.175 76.745 ;
        RECT 143.345 76.805 143.605 77.065 ;
        RECT 143.345 76.485 143.605 76.745 ;
        RECT 143.775 76.805 144.035 77.065 ;
        RECT 143.775 76.485 144.035 76.745 ;
        RECT 144.205 76.805 144.465 77.065 ;
        RECT 144.205 76.485 144.465 76.745 ;
        RECT 144.635 76.805 144.895 77.065 ;
        RECT 144.635 76.485 144.895 76.745 ;
        RECT 145.065 76.805 145.325 77.065 ;
        RECT 145.065 76.485 145.325 76.745 ;
        RECT 145.495 76.805 145.755 77.065 ;
        RECT 145.495 76.485 145.755 76.745 ;
        RECT 145.925 76.805 146.185 77.065 ;
        RECT 145.925 76.485 146.185 76.745 ;
        RECT 146.355 76.805 146.615 77.065 ;
        RECT 146.355 76.485 146.615 76.745 ;
        RECT 146.985 76.805 147.245 77.065 ;
        RECT 146.985 76.485 147.245 76.745 ;
        RECT 43.505 74.715 43.765 74.975 ;
        RECT 43.825 74.715 44.085 74.975 ;
        RECT 44.145 74.715 44.405 74.975 ;
        RECT 44.465 74.715 44.725 74.975 ;
        RECT 44.785 74.715 45.045 74.975 ;
        RECT 45.105 74.715 45.365 74.975 ;
        RECT 45.425 74.715 45.685 74.975 ;
        RECT 45.745 74.715 46.005 74.975 ;
        RECT 46.065 74.715 46.325 74.975 ;
        RECT 46.385 74.715 46.645 74.975 ;
        RECT 46.705 74.715 46.965 74.975 ;
        RECT 47.025 74.715 47.285 74.975 ;
        RECT 47.345 74.715 47.605 74.975 ;
        RECT 47.665 74.715 47.925 74.975 ;
        RECT 47.985 74.715 48.245 74.975 ;
        RECT 48.305 74.715 48.565 74.975 ;
        RECT 48.625 74.715 48.885 74.975 ;
        RECT 48.945 74.715 49.205 74.975 ;
        RECT 49.265 74.715 49.525 74.975 ;
        RECT 49.585 74.715 49.845 74.975 ;
        RECT 49.905 74.715 50.165 74.975 ;
        RECT 50.225 74.715 50.485 74.975 ;
        RECT 50.545 74.715 50.805 74.975 ;
        RECT 50.865 74.715 51.125 74.975 ;
        RECT 51.185 74.715 51.445 74.975 ;
        RECT 51.505 74.715 51.765 74.975 ;
        RECT 51.825 74.715 52.085 74.975 ;
        RECT 52.145 74.715 52.405 74.975 ;
        RECT 52.465 74.715 52.725 74.975 ;
        RECT 52.785 74.715 53.045 74.975 ;
        RECT 53.105 74.715 53.365 74.975 ;
        RECT 53.425 74.715 53.685 74.975 ;
        RECT 53.745 74.715 54.005 74.975 ;
        RECT 54.065 74.715 54.325 74.975 ;
        RECT 54.385 74.715 54.645 74.975 ;
        RECT 54.705 74.715 54.965 74.975 ;
        RECT 55.025 74.715 55.285 74.975 ;
        RECT 55.345 74.715 55.605 74.975 ;
        RECT 55.665 74.715 55.925 74.975 ;
        RECT 55.985 74.715 56.245 74.975 ;
        RECT 56.305 74.715 56.565 74.975 ;
        RECT 56.625 74.715 56.885 74.975 ;
        RECT 56.945 74.715 57.205 74.975 ;
        RECT 57.265 74.715 57.525 74.975 ;
        RECT 57.585 74.715 57.845 74.975 ;
        RECT 57.905 74.715 58.165 74.975 ;
        RECT 58.225 74.715 58.485 74.975 ;
        RECT 58.545 74.715 58.805 74.975 ;
        RECT 58.865 74.715 59.125 74.975 ;
        RECT 59.185 74.715 59.445 74.975 ;
        RECT 59.505 74.715 59.765 74.975 ;
        RECT 59.825 74.715 60.085 74.975 ;
        RECT 60.145 74.715 60.405 74.975 ;
        RECT 60.465 74.715 60.725 74.975 ;
        RECT 60.785 74.715 61.045 74.975 ;
        RECT 61.105 74.715 61.365 74.975 ;
        RECT 61.425 74.715 61.685 74.975 ;
        RECT 61.745 74.715 62.005 74.975 ;
        RECT 62.065 74.715 62.325 74.975 ;
        RECT 62.385 74.715 62.645 74.975 ;
        RECT 62.705 74.715 62.965 74.975 ;
        RECT 63.025 74.715 63.285 74.975 ;
        RECT 63.345 74.715 63.605 74.975 ;
        RECT 63.665 74.715 63.925 74.975 ;
        RECT 63.985 74.715 64.245 74.975 ;
        RECT 64.305 74.715 64.565 74.975 ;
        RECT 64.625 74.715 64.885 74.975 ;
        RECT 64.945 74.715 65.205 74.975 ;
        RECT 65.265 74.715 65.525 74.975 ;
        RECT 65.585 74.715 65.845 74.975 ;
        RECT 65.905 74.715 66.165 74.975 ;
        RECT 66.225 74.715 66.485 74.975 ;
        RECT 66.545 74.715 66.805 74.975 ;
        RECT 66.865 74.715 67.125 74.975 ;
        RECT 67.185 74.715 67.445 74.975 ;
        RECT 67.505 74.715 67.765 74.975 ;
        RECT 67.825 74.715 68.085 74.975 ;
        RECT 68.145 74.715 68.405 74.975 ;
        RECT 68.465 74.715 68.725 74.975 ;
        RECT 68.785 74.715 69.045 74.975 ;
        RECT 69.105 74.715 69.365 74.975 ;
        RECT 69.425 74.715 69.685 74.975 ;
        RECT 69.745 74.715 70.005 74.975 ;
        RECT 70.065 74.715 70.325 74.975 ;
        RECT 70.385 74.715 70.645 74.975 ;
        RECT 70.705 74.715 70.965 74.975 ;
        RECT 123.980 74.715 124.240 74.975 ;
        RECT 124.300 74.715 124.560 74.975 ;
        RECT 124.620 74.715 124.880 74.975 ;
        RECT 42.725 74.190 42.985 74.450 ;
        RECT 42.725 73.870 42.985 74.130 ;
        RECT 43.355 74.190 43.615 74.450 ;
        RECT 43.355 73.870 43.615 74.130 ;
        RECT 45.635 74.190 45.895 74.450 ;
        RECT 45.635 73.870 45.895 74.130 ;
        RECT 47.915 74.190 48.175 74.450 ;
        RECT 47.915 73.870 48.175 74.130 ;
        RECT 50.195 74.190 50.455 74.450 ;
        RECT 50.195 73.870 50.455 74.130 ;
        RECT 52.475 74.190 52.735 74.450 ;
        RECT 52.475 73.870 52.735 74.130 ;
        RECT 54.755 74.190 55.015 74.450 ;
        RECT 54.755 73.870 55.015 74.130 ;
        RECT 57.035 74.190 57.295 74.450 ;
        RECT 57.035 73.870 57.295 74.130 ;
        RECT 59.315 74.190 59.575 74.450 ;
        RECT 59.315 73.870 59.575 74.130 ;
        RECT 61.595 74.190 61.855 74.450 ;
        RECT 61.595 73.870 61.855 74.130 ;
        RECT 63.875 74.190 64.135 74.450 ;
        RECT 63.875 73.870 64.135 74.130 ;
        RECT 66.155 74.190 66.415 74.450 ;
        RECT 66.155 73.870 66.415 74.130 ;
        RECT 68.435 74.190 68.695 74.450 ;
        RECT 68.435 73.870 68.695 74.130 ;
        RECT 70.715 74.190 70.975 74.450 ;
        RECT 70.715 73.870 70.975 74.130 ;
        RECT 72.995 74.190 73.255 74.450 ;
        RECT 72.995 73.870 73.255 74.130 ;
        RECT 75.275 74.190 75.535 74.450 ;
        RECT 75.275 73.870 75.535 74.130 ;
        RECT 77.555 74.190 77.815 74.450 ;
        RECT 77.555 73.870 77.815 74.130 ;
        RECT 79.835 74.190 80.095 74.450 ;
        RECT 79.835 73.870 80.095 74.130 ;
        RECT 82.115 74.190 82.375 74.450 ;
        RECT 82.115 73.870 82.375 74.130 ;
        RECT 84.395 74.190 84.655 74.450 ;
        RECT 84.395 73.870 84.655 74.130 ;
        RECT 86.675 74.190 86.935 74.450 ;
        RECT 86.675 73.870 86.935 74.130 ;
        RECT 88.955 74.190 89.215 74.450 ;
        RECT 88.955 73.870 89.215 74.130 ;
        RECT 91.235 74.190 91.495 74.450 ;
        RECT 91.235 73.870 91.495 74.130 ;
        RECT 93.515 74.190 93.775 74.450 ;
        RECT 93.515 73.870 93.775 74.130 ;
        RECT 95.795 74.190 96.055 74.450 ;
        RECT 95.795 73.870 96.055 74.130 ;
        RECT 98.075 74.190 98.335 74.450 ;
        RECT 98.075 73.870 98.335 74.130 ;
        RECT 100.355 74.190 100.615 74.450 ;
        RECT 100.355 73.870 100.615 74.130 ;
        RECT 102.635 74.190 102.895 74.450 ;
        RECT 102.635 73.870 102.895 74.130 ;
        RECT 104.915 74.190 105.175 74.450 ;
        RECT 104.915 73.870 105.175 74.130 ;
        RECT 107.195 74.190 107.455 74.450 ;
        RECT 107.195 73.870 107.455 74.130 ;
        RECT 109.475 74.190 109.735 74.450 ;
        RECT 109.475 73.870 109.735 74.130 ;
        RECT 111.755 74.190 112.015 74.450 ;
        RECT 111.755 73.870 112.015 74.130 ;
        RECT 114.035 74.190 114.295 74.450 ;
        RECT 114.035 73.870 114.295 74.130 ;
        RECT 116.315 74.190 116.575 74.450 ;
        RECT 116.315 73.870 116.575 74.130 ;
        RECT 118.595 74.190 118.855 74.450 ;
        RECT 118.595 73.870 118.855 74.130 ;
        RECT 120.875 74.190 121.135 74.450 ;
        RECT 120.875 73.870 121.135 74.130 ;
        RECT 123.155 74.190 123.415 74.450 ;
        RECT 123.155 73.870 123.415 74.130 ;
        RECT 125.435 74.190 125.695 74.450 ;
        RECT 125.435 73.870 125.695 74.130 ;
        RECT 127.715 74.190 127.975 74.450 ;
        RECT 127.715 73.870 127.975 74.130 ;
        RECT 129.995 74.190 130.255 74.450 ;
        RECT 129.995 73.870 130.255 74.130 ;
        RECT 130.625 74.190 130.885 74.450 ;
        RECT 130.625 73.870 130.885 74.130 ;
        RECT 123.980 73.345 124.240 73.605 ;
        RECT 124.300 73.345 124.560 73.605 ;
        RECT 124.620 73.345 124.880 73.605 ;
        RECT 137.660 74.080 137.920 74.340 ;
        RECT 137.980 74.080 138.240 74.340 ;
        RECT 138.300 74.080 138.560 74.340 ;
        RECT 138.615 73.535 138.875 73.795 ;
        RECT 138.615 73.215 138.875 73.475 ;
        RECT 139.045 73.535 139.305 73.795 ;
        RECT 139.045 73.215 139.305 73.475 ;
        RECT 139.475 73.535 139.735 73.795 ;
        RECT 139.475 73.215 139.735 73.475 ;
        RECT 139.905 73.535 140.165 73.795 ;
        RECT 139.905 73.215 140.165 73.475 ;
        RECT 140.335 73.535 140.595 73.795 ;
        RECT 140.335 73.215 140.595 73.475 ;
        RECT 93.260 71.390 93.520 71.650 ;
        RECT 93.580 71.390 93.840 71.650 ;
        RECT 93.900 71.390 94.160 71.650 ;
        RECT 93.155 70.855 93.415 71.115 ;
        RECT 93.155 70.535 93.415 70.795 ;
        RECT 93.155 70.215 93.415 70.475 ;
        RECT 94.015 70.855 94.275 71.115 ;
        RECT 94.015 70.535 94.275 70.795 ;
        RECT 94.015 70.215 94.275 70.475 ;
        RECT 127.460 71.390 127.720 71.650 ;
        RECT 127.780 71.390 128.040 71.650 ;
        RECT 128.100 71.390 128.360 71.650 ;
        RECT 127.355 70.855 127.615 71.115 ;
        RECT 127.355 70.535 127.615 70.795 ;
        RECT 127.355 70.215 127.615 70.475 ;
        RECT 128.215 70.855 128.475 71.115 ;
        RECT 128.215 70.535 128.475 70.795 ;
        RECT 128.215 70.215 128.475 70.475 ;
        RECT 137.670 71.365 137.930 71.625 ;
        RECT 137.990 71.365 138.250 71.625 ;
        RECT 137.085 70.820 137.345 71.080 ;
        RECT 137.085 70.500 137.345 70.760 ;
        RECT 137.755 70.820 138.015 71.080 ;
        RECT 137.755 70.500 138.015 70.760 ;
        RECT 138.185 70.820 138.445 71.080 ;
        RECT 138.185 70.500 138.445 70.760 ;
        RECT 138.615 70.820 138.875 71.080 ;
        RECT 138.615 70.500 138.875 70.760 ;
        RECT 139.030 70.820 139.290 71.080 ;
        RECT 139.030 70.500 139.290 70.760 ;
        RECT 139.475 70.820 139.735 71.080 ;
        RECT 139.475 70.500 139.735 70.760 ;
        RECT 139.890 70.820 140.150 71.080 ;
        RECT 139.890 70.500 140.150 70.760 ;
        RECT 140.335 70.820 140.595 71.080 ;
        RECT 140.335 70.500 140.595 70.760 ;
        RECT 140.765 70.820 141.025 71.080 ;
        RECT 140.765 70.500 141.025 70.760 ;
        RECT 141.195 70.820 141.455 71.080 ;
        RECT 141.195 70.500 141.455 70.760 ;
        RECT 145.970 74.080 146.230 74.340 ;
        RECT 146.290 74.080 146.550 74.340 ;
        RECT 143.865 73.535 144.125 73.795 ;
        RECT 143.865 73.215 144.125 73.475 ;
        RECT 144.295 73.535 144.555 73.795 ;
        RECT 144.295 73.215 144.555 73.475 ;
        RECT 144.725 73.535 144.985 73.795 ;
        RECT 144.725 73.215 144.985 73.475 ;
        RECT 145.155 73.535 145.415 73.795 ;
        RECT 145.155 73.215 145.415 73.475 ;
        RECT 145.585 73.535 145.845 73.795 ;
        RECT 145.585 73.215 145.845 73.475 ;
        RECT 143.030 71.475 143.290 71.735 ;
        RECT 143.350 71.475 143.610 71.735 ;
        RECT 143.670 71.475 143.930 71.735 ;
        RECT 143.005 70.820 143.265 71.080 ;
        RECT 143.005 70.500 143.265 70.760 ;
        RECT 143.435 70.820 143.695 71.080 ;
        RECT 143.435 70.500 143.695 70.760 ;
        RECT 143.865 70.820 144.125 71.080 ;
        RECT 143.865 70.500 144.125 70.760 ;
        RECT 144.280 70.820 144.540 71.080 ;
        RECT 144.280 70.500 144.540 70.760 ;
        RECT 144.725 70.820 144.985 71.080 ;
        RECT 144.725 70.500 144.985 70.760 ;
        RECT 145.140 70.820 145.400 71.080 ;
        RECT 145.140 70.500 145.400 70.760 ;
        RECT 145.585 70.820 145.845 71.080 ;
        RECT 145.585 70.500 145.845 70.760 ;
        RECT 146.015 70.820 146.275 71.080 ;
        RECT 146.015 70.500 146.275 70.760 ;
        RECT 146.445 70.820 146.705 71.080 ;
        RECT 146.445 70.500 146.705 70.760 ;
        RECT 147.075 70.820 147.335 71.080 ;
        RECT 147.075 70.500 147.335 70.760 ;
        RECT 90.770 67.275 91.030 67.535 ;
        RECT 90.770 66.955 91.030 67.215 ;
        RECT 91.200 67.275 91.460 67.535 ;
        RECT 91.200 66.955 91.460 67.215 ;
        RECT 91.630 67.275 91.890 67.535 ;
        RECT 91.630 66.955 91.890 67.215 ;
        RECT 90.315 66.410 90.575 66.670 ;
        RECT 90.635 66.410 90.895 66.670 ;
        RECT 96.865 67.820 97.125 68.080 ;
        RECT 97.185 67.820 97.445 68.080 ;
        RECT 95.440 67.275 95.700 67.535 ;
        RECT 95.440 66.955 95.700 67.215 ;
        RECT 95.870 67.275 96.130 67.535 ;
        RECT 95.870 66.955 96.130 67.215 ;
        RECT 96.300 67.275 96.560 67.535 ;
        RECT 96.300 66.955 96.560 67.215 ;
        RECT 124.970 67.275 125.230 67.535 ;
        RECT 124.970 66.955 125.230 67.215 ;
        RECT 125.400 67.275 125.660 67.535 ;
        RECT 125.400 66.955 125.660 67.215 ;
        RECT 125.830 67.275 126.090 67.535 ;
        RECT 125.830 66.955 126.090 67.215 ;
        RECT 124.515 66.410 124.775 66.670 ;
        RECT 124.835 66.410 125.095 66.670 ;
        RECT 131.065 67.820 131.325 68.080 ;
        RECT 131.385 67.820 131.645 68.080 ;
        RECT 129.640 67.275 129.900 67.535 ;
        RECT 129.640 66.955 129.900 67.215 ;
        RECT 130.070 67.275 130.330 67.535 ;
        RECT 130.070 66.955 130.330 67.215 ;
        RECT 130.500 67.275 130.760 67.535 ;
        RECT 130.500 66.955 130.760 67.215 ;
        RECT 132.030 67.125 132.290 67.385 ;
        RECT 132.030 66.805 132.290 67.065 ;
        RECT 136.805 67.125 137.065 67.385 ;
        RECT 136.805 66.805 137.065 67.065 ;
        RECT 137.475 67.125 137.735 67.385 ;
        RECT 137.475 66.805 137.735 67.065 ;
        RECT 139.755 67.125 140.015 67.385 ;
        RECT 139.755 66.805 140.015 67.065 ;
        RECT 142.035 67.125 142.295 67.385 ;
        RECT 142.035 66.805 142.295 67.065 ;
        RECT 144.315 67.125 144.575 67.385 ;
        RECT 144.315 66.805 144.575 67.065 ;
        RECT 146.595 67.125 146.855 67.385 ;
        RECT 146.595 66.805 146.855 67.065 ;
        RECT 147.265 67.125 147.525 67.385 ;
        RECT 147.265 66.805 147.525 67.065 ;
        RECT 137.960 66.260 138.220 66.520 ;
        RECT 138.280 66.260 138.540 66.520 ;
        RECT 138.600 66.260 138.860 66.520 ;
        RECT 35.495 64.215 35.755 64.475 ;
        RECT 33.535 63.735 33.795 63.995 ;
        RECT 33.535 63.415 33.795 63.675 ;
        RECT 33.535 63.095 33.795 63.355 ;
        RECT 34.205 63.735 34.465 63.995 ;
        RECT 34.205 63.415 34.465 63.675 ;
        RECT 34.205 63.095 34.465 63.355 ;
        RECT 34.635 63.735 34.895 63.995 ;
        RECT 34.635 63.415 34.895 63.675 ;
        RECT 34.635 63.095 34.895 63.355 ;
        RECT 35.065 63.735 35.325 63.995 ;
        RECT 35.065 63.415 35.325 63.675 ;
        RECT 35.065 63.095 35.325 63.355 ;
        RECT 35.495 63.895 35.755 64.155 ;
        RECT 36.355 64.215 36.615 64.475 ;
        RECT 35.495 63.575 35.755 63.835 ;
        RECT 35.495 63.255 35.755 63.515 ;
        RECT 35.495 62.935 35.755 63.195 ;
        RECT 35.925 63.735 36.185 63.995 ;
        RECT 35.925 63.415 36.185 63.675 ;
        RECT 35.925 63.095 36.185 63.355 ;
        RECT 36.355 63.895 36.615 64.155 ;
        RECT 36.355 63.575 36.615 63.835 ;
        RECT 36.355 63.255 36.615 63.515 ;
        RECT 35.495 62.615 35.755 62.875 ;
        RECT 36.355 62.935 36.615 63.195 ;
        RECT 36.785 63.735 37.045 63.995 ;
        RECT 36.785 63.415 37.045 63.675 ;
        RECT 36.785 63.095 37.045 63.355 ;
        RECT 37.215 63.735 37.475 63.995 ;
        RECT 37.215 63.415 37.475 63.675 ;
        RECT 37.215 63.095 37.475 63.355 ;
        RECT 37.645 63.735 37.905 63.995 ;
        RECT 37.645 63.415 37.905 63.675 ;
        RECT 37.645 63.095 37.905 63.355 ;
        RECT 38.315 63.735 38.575 63.995 ;
        RECT 38.315 63.415 38.575 63.675 ;
        RECT 38.315 63.095 38.575 63.355 ;
        RECT 36.355 62.615 36.615 62.875 ;
        RECT 42.685 63.725 42.945 63.985 ;
        RECT 42.685 63.405 42.945 63.665 ;
        RECT 43.355 63.725 43.615 63.985 ;
        RECT 43.355 63.405 43.615 63.665 ;
        RECT 45.635 63.725 45.895 63.985 ;
        RECT 45.635 63.405 45.895 63.665 ;
        RECT 47.915 63.725 48.175 63.985 ;
        RECT 47.915 63.405 48.175 63.665 ;
        RECT 50.195 63.725 50.455 63.985 ;
        RECT 50.195 63.405 50.455 63.665 ;
        RECT 52.475 63.725 52.735 63.985 ;
        RECT 52.475 63.405 52.735 63.665 ;
        RECT 54.755 63.725 55.015 63.985 ;
        RECT 54.755 63.405 55.015 63.665 ;
        RECT 57.035 63.725 57.295 63.985 ;
        RECT 57.035 63.405 57.295 63.665 ;
        RECT 59.315 63.725 59.575 63.985 ;
        RECT 59.315 63.405 59.575 63.665 ;
        RECT 61.595 63.725 61.855 63.985 ;
        RECT 61.595 63.405 61.855 63.665 ;
        RECT 63.875 63.725 64.135 63.985 ;
        RECT 63.875 63.405 64.135 63.665 ;
        RECT 66.155 63.725 66.415 63.985 ;
        RECT 66.155 63.405 66.415 63.665 ;
        RECT 68.435 63.725 68.695 63.985 ;
        RECT 68.435 63.405 68.695 63.665 ;
        RECT 70.715 63.725 70.975 63.985 ;
        RECT 70.715 63.405 70.975 63.665 ;
        RECT 72.995 63.725 73.255 63.985 ;
        RECT 72.995 63.405 73.255 63.665 ;
        RECT 75.275 63.725 75.535 63.985 ;
        RECT 75.275 63.405 75.535 63.665 ;
        RECT 77.555 63.725 77.815 63.985 ;
        RECT 77.555 63.405 77.815 63.665 ;
        RECT 79.835 63.725 80.095 63.985 ;
        RECT 79.835 63.405 80.095 63.665 ;
        RECT 82.115 63.725 82.375 63.985 ;
        RECT 82.115 63.405 82.375 63.665 ;
        RECT 84.395 63.725 84.655 63.985 ;
        RECT 84.395 63.405 84.655 63.665 ;
        RECT 86.675 63.725 86.935 63.985 ;
        RECT 86.675 63.405 86.935 63.665 ;
        RECT 88.955 63.725 89.215 63.985 ;
        RECT 88.955 63.405 89.215 63.665 ;
        RECT 91.235 63.725 91.495 63.985 ;
        RECT 91.235 63.405 91.495 63.665 ;
        RECT 93.515 63.725 93.775 63.985 ;
        RECT 93.515 63.405 93.775 63.665 ;
        RECT 95.795 63.725 96.055 63.985 ;
        RECT 95.795 63.405 96.055 63.665 ;
        RECT 98.075 63.725 98.335 63.985 ;
        RECT 98.075 63.405 98.335 63.665 ;
        RECT 100.355 63.725 100.615 63.985 ;
        RECT 100.355 63.405 100.615 63.665 ;
        RECT 102.635 63.725 102.895 63.985 ;
        RECT 102.635 63.405 102.895 63.665 ;
        RECT 104.915 63.725 105.175 63.985 ;
        RECT 104.915 63.405 105.175 63.665 ;
        RECT 107.195 63.725 107.455 63.985 ;
        RECT 107.195 63.405 107.455 63.665 ;
        RECT 109.475 63.725 109.735 63.985 ;
        RECT 109.475 63.405 109.735 63.665 ;
        RECT 111.755 63.725 112.015 63.985 ;
        RECT 111.755 63.405 112.015 63.665 ;
        RECT 114.035 63.725 114.295 63.985 ;
        RECT 114.035 63.405 114.295 63.665 ;
        RECT 116.315 63.725 116.575 63.985 ;
        RECT 116.315 63.405 116.575 63.665 ;
        RECT 118.595 63.725 118.855 63.985 ;
        RECT 118.595 63.405 118.855 63.665 ;
        RECT 120.875 63.725 121.135 63.985 ;
        RECT 120.875 63.405 121.135 63.665 ;
        RECT 123.155 63.725 123.415 63.985 ;
        RECT 123.155 63.405 123.415 63.665 ;
        RECT 125.435 63.725 125.695 63.985 ;
        RECT 125.435 63.405 125.695 63.665 ;
        RECT 127.715 63.725 127.975 63.985 ;
        RECT 127.715 63.405 127.975 63.665 ;
        RECT 129.995 63.725 130.255 63.985 ;
        RECT 129.995 63.405 130.255 63.665 ;
        RECT 132.275 63.725 132.535 63.985 ;
        RECT 132.275 63.405 132.535 63.665 ;
        RECT 134.555 63.725 134.815 63.985 ;
        RECT 134.555 63.405 134.815 63.665 ;
        RECT 136.835 63.725 137.095 63.985 ;
        RECT 136.835 63.405 137.095 63.665 ;
        RECT 139.115 63.725 139.375 63.985 ;
        RECT 139.115 63.405 139.375 63.665 ;
        RECT 141.395 63.725 141.655 63.985 ;
        RECT 141.395 63.405 141.655 63.665 ;
        RECT 143.675 63.725 143.935 63.985 ;
        RECT 143.675 63.405 143.935 63.665 ;
        RECT 144.345 63.725 144.605 63.985 ;
        RECT 144.345 63.405 144.605 63.665 ;
        RECT 107.895 62.880 108.155 63.140 ;
        RECT 108.215 62.880 108.475 63.140 ;
        RECT 108.535 62.880 108.795 63.140 ;
        RECT 108.855 62.880 109.115 63.140 ;
        RECT 137.650 62.880 137.910 63.140 ;
        RECT 137.970 62.880 138.230 63.140 ;
        RECT 138.290 62.880 138.550 63.140 ;
        RECT 42.685 62.355 42.945 62.615 ;
        RECT 42.685 62.035 42.945 62.295 ;
        RECT 43.355 62.355 43.615 62.615 ;
        RECT 43.355 62.035 43.615 62.295 ;
        RECT 45.635 62.355 45.895 62.615 ;
        RECT 45.635 62.035 45.895 62.295 ;
        RECT 47.915 62.355 48.175 62.615 ;
        RECT 47.915 62.035 48.175 62.295 ;
        RECT 50.195 62.355 50.455 62.615 ;
        RECT 50.195 62.035 50.455 62.295 ;
        RECT 52.475 62.355 52.735 62.615 ;
        RECT 52.475 62.035 52.735 62.295 ;
        RECT 54.755 62.355 55.015 62.615 ;
        RECT 54.755 62.035 55.015 62.295 ;
        RECT 57.035 62.355 57.295 62.615 ;
        RECT 57.035 62.035 57.295 62.295 ;
        RECT 59.315 62.355 59.575 62.615 ;
        RECT 59.315 62.035 59.575 62.295 ;
        RECT 61.595 62.355 61.855 62.615 ;
        RECT 61.595 62.035 61.855 62.295 ;
        RECT 63.875 62.355 64.135 62.615 ;
        RECT 63.875 62.035 64.135 62.295 ;
        RECT 66.155 62.355 66.415 62.615 ;
        RECT 66.155 62.035 66.415 62.295 ;
        RECT 68.435 62.355 68.695 62.615 ;
        RECT 68.435 62.035 68.695 62.295 ;
        RECT 70.715 62.355 70.975 62.615 ;
        RECT 70.715 62.035 70.975 62.295 ;
        RECT 72.995 62.355 73.255 62.615 ;
        RECT 72.995 62.035 73.255 62.295 ;
        RECT 75.275 62.355 75.535 62.615 ;
        RECT 75.275 62.035 75.535 62.295 ;
        RECT 77.555 62.355 77.815 62.615 ;
        RECT 77.555 62.035 77.815 62.295 ;
        RECT 79.835 62.355 80.095 62.615 ;
        RECT 79.835 62.035 80.095 62.295 ;
        RECT 82.115 62.355 82.375 62.615 ;
        RECT 82.115 62.035 82.375 62.295 ;
        RECT 84.395 62.355 84.655 62.615 ;
        RECT 84.395 62.035 84.655 62.295 ;
        RECT 86.675 62.355 86.935 62.615 ;
        RECT 86.675 62.035 86.935 62.295 ;
        RECT 88.955 62.355 89.215 62.615 ;
        RECT 88.955 62.035 89.215 62.295 ;
        RECT 91.235 62.355 91.495 62.615 ;
        RECT 91.235 62.035 91.495 62.295 ;
        RECT 93.515 62.355 93.775 62.615 ;
        RECT 93.515 62.035 93.775 62.295 ;
        RECT 95.795 62.355 96.055 62.615 ;
        RECT 95.795 62.035 96.055 62.295 ;
        RECT 98.075 62.355 98.335 62.615 ;
        RECT 98.075 62.035 98.335 62.295 ;
        RECT 100.355 62.355 100.615 62.615 ;
        RECT 100.355 62.035 100.615 62.295 ;
        RECT 102.635 62.355 102.895 62.615 ;
        RECT 102.635 62.035 102.895 62.295 ;
        RECT 104.915 62.355 105.175 62.615 ;
        RECT 104.915 62.035 105.175 62.295 ;
        RECT 107.195 62.355 107.455 62.615 ;
        RECT 107.195 62.035 107.455 62.295 ;
        RECT 109.475 62.355 109.735 62.615 ;
        RECT 109.475 62.035 109.735 62.295 ;
        RECT 111.755 62.355 112.015 62.615 ;
        RECT 111.755 62.035 112.015 62.295 ;
        RECT 114.035 62.355 114.295 62.615 ;
        RECT 114.035 62.035 114.295 62.295 ;
        RECT 116.315 62.355 116.575 62.615 ;
        RECT 116.315 62.035 116.575 62.295 ;
        RECT 118.595 62.355 118.855 62.615 ;
        RECT 118.595 62.035 118.855 62.295 ;
        RECT 120.875 62.355 121.135 62.615 ;
        RECT 120.875 62.035 121.135 62.295 ;
        RECT 123.155 62.355 123.415 62.615 ;
        RECT 123.155 62.035 123.415 62.295 ;
        RECT 125.435 62.355 125.695 62.615 ;
        RECT 125.435 62.035 125.695 62.295 ;
        RECT 127.715 62.355 127.975 62.615 ;
        RECT 127.715 62.035 127.975 62.295 ;
        RECT 129.995 62.355 130.255 62.615 ;
        RECT 129.995 62.035 130.255 62.295 ;
        RECT 132.275 62.355 132.535 62.615 ;
        RECT 132.275 62.035 132.535 62.295 ;
        RECT 134.555 62.355 134.815 62.615 ;
        RECT 134.555 62.035 134.815 62.295 ;
        RECT 136.835 62.355 137.095 62.615 ;
        RECT 136.835 62.035 137.095 62.295 ;
        RECT 139.115 62.355 139.375 62.615 ;
        RECT 139.115 62.035 139.375 62.295 ;
        RECT 141.395 62.355 141.655 62.615 ;
        RECT 141.395 62.035 141.655 62.295 ;
        RECT 143.675 62.355 143.935 62.615 ;
        RECT 143.675 62.035 143.935 62.295 ;
        RECT 144.345 62.355 144.605 62.615 ;
        RECT 144.345 62.035 144.605 62.295 ;
        RECT 34.300 61.240 34.560 61.500 ;
        RECT 34.620 61.240 34.880 61.500 ;
        RECT 33.535 59.885 33.795 60.145 ;
        RECT 33.535 59.565 33.795 59.825 ;
        RECT 33.535 59.245 33.795 59.505 ;
        RECT 34.205 59.885 34.465 60.145 ;
        RECT 34.205 59.565 34.465 59.825 ;
        RECT 34.205 59.245 34.465 59.505 ;
        RECT 34.635 59.885 34.895 60.145 ;
        RECT 34.635 59.565 34.895 59.825 ;
        RECT 34.635 59.245 34.895 59.505 ;
        RECT 35.065 59.885 35.325 60.145 ;
        RECT 35.065 59.565 35.325 59.825 ;
        RECT 35.065 59.245 35.325 59.505 ;
        RECT 35.495 59.885 35.755 60.145 ;
        RECT 35.495 59.565 35.755 59.825 ;
        RECT 35.495 59.245 35.755 59.505 ;
        RECT 35.925 59.885 36.185 60.145 ;
        RECT 35.925 59.565 36.185 59.825 ;
        RECT 35.925 59.245 36.185 59.505 ;
        RECT 36.355 59.885 36.615 60.145 ;
        RECT 36.355 59.565 36.615 59.825 ;
        RECT 36.355 59.245 36.615 59.505 ;
        RECT 36.785 59.885 37.045 60.145 ;
        RECT 36.785 59.565 37.045 59.825 ;
        RECT 36.785 59.245 37.045 59.505 ;
        RECT 37.215 59.885 37.475 60.145 ;
        RECT 37.215 59.565 37.475 59.825 ;
        RECT 37.215 59.245 37.475 59.505 ;
        RECT 37.645 59.885 37.905 60.145 ;
        RECT 37.645 59.565 37.905 59.825 ;
        RECT 37.645 59.245 37.905 59.505 ;
        RECT 38.315 59.885 38.575 60.145 ;
        RECT 38.315 59.565 38.575 59.825 ;
        RECT 42.685 60.985 42.945 61.245 ;
        RECT 42.685 60.665 42.945 60.925 ;
        RECT 43.355 60.985 43.615 61.245 ;
        RECT 43.355 60.665 43.615 60.925 ;
        RECT 45.635 60.985 45.895 61.245 ;
        RECT 45.635 60.665 45.895 60.925 ;
        RECT 47.915 60.985 48.175 61.245 ;
        RECT 47.915 60.665 48.175 60.925 ;
        RECT 50.195 60.985 50.455 61.245 ;
        RECT 50.195 60.665 50.455 60.925 ;
        RECT 52.475 60.985 52.735 61.245 ;
        RECT 52.475 60.665 52.735 60.925 ;
        RECT 54.755 60.985 55.015 61.245 ;
        RECT 54.755 60.665 55.015 60.925 ;
        RECT 57.035 60.985 57.295 61.245 ;
        RECT 57.035 60.665 57.295 60.925 ;
        RECT 59.315 60.985 59.575 61.245 ;
        RECT 59.315 60.665 59.575 60.925 ;
        RECT 61.595 60.985 61.855 61.245 ;
        RECT 61.595 60.665 61.855 60.925 ;
        RECT 63.875 60.985 64.135 61.245 ;
        RECT 63.875 60.665 64.135 60.925 ;
        RECT 66.155 60.985 66.415 61.245 ;
        RECT 66.155 60.665 66.415 60.925 ;
        RECT 68.435 60.985 68.695 61.245 ;
        RECT 68.435 60.665 68.695 60.925 ;
        RECT 70.715 60.985 70.975 61.245 ;
        RECT 70.715 60.665 70.975 60.925 ;
        RECT 72.995 60.985 73.255 61.245 ;
        RECT 72.995 60.665 73.255 60.925 ;
        RECT 75.275 60.985 75.535 61.245 ;
        RECT 75.275 60.665 75.535 60.925 ;
        RECT 77.555 60.985 77.815 61.245 ;
        RECT 77.555 60.665 77.815 60.925 ;
        RECT 79.835 60.985 80.095 61.245 ;
        RECT 79.835 60.665 80.095 60.925 ;
        RECT 82.115 60.985 82.375 61.245 ;
        RECT 82.115 60.665 82.375 60.925 ;
        RECT 84.395 60.985 84.655 61.245 ;
        RECT 84.395 60.665 84.655 60.925 ;
        RECT 86.675 60.985 86.935 61.245 ;
        RECT 86.675 60.665 86.935 60.925 ;
        RECT 88.955 60.985 89.215 61.245 ;
        RECT 88.955 60.665 89.215 60.925 ;
        RECT 91.235 60.985 91.495 61.245 ;
        RECT 91.235 60.665 91.495 60.925 ;
        RECT 93.515 60.985 93.775 61.245 ;
        RECT 93.515 60.665 93.775 60.925 ;
        RECT 95.795 60.985 96.055 61.245 ;
        RECT 95.795 60.665 96.055 60.925 ;
        RECT 98.075 60.985 98.335 61.245 ;
        RECT 98.075 60.665 98.335 60.925 ;
        RECT 100.355 60.985 100.615 61.245 ;
        RECT 100.355 60.665 100.615 60.925 ;
        RECT 102.635 60.985 102.895 61.245 ;
        RECT 102.635 60.665 102.895 60.925 ;
        RECT 104.915 60.985 105.175 61.245 ;
        RECT 104.915 60.665 105.175 60.925 ;
        RECT 107.195 60.985 107.455 61.245 ;
        RECT 107.195 60.665 107.455 60.925 ;
        RECT 109.475 60.985 109.735 61.245 ;
        RECT 109.475 60.665 109.735 60.925 ;
        RECT 111.755 60.985 112.015 61.245 ;
        RECT 111.755 60.665 112.015 60.925 ;
        RECT 114.035 60.985 114.295 61.245 ;
        RECT 114.035 60.665 114.295 60.925 ;
        RECT 116.315 60.985 116.575 61.245 ;
        RECT 116.315 60.665 116.575 60.925 ;
        RECT 118.595 60.985 118.855 61.245 ;
        RECT 118.595 60.665 118.855 60.925 ;
        RECT 120.875 60.985 121.135 61.245 ;
        RECT 120.875 60.665 121.135 60.925 ;
        RECT 123.155 60.985 123.415 61.245 ;
        RECT 123.155 60.665 123.415 60.925 ;
        RECT 125.435 60.985 125.695 61.245 ;
        RECT 125.435 60.665 125.695 60.925 ;
        RECT 127.715 60.985 127.975 61.245 ;
        RECT 127.715 60.665 127.975 60.925 ;
        RECT 129.995 60.985 130.255 61.245 ;
        RECT 129.995 60.665 130.255 60.925 ;
        RECT 132.275 60.985 132.535 61.245 ;
        RECT 132.275 60.665 132.535 60.925 ;
        RECT 134.555 60.985 134.815 61.245 ;
        RECT 134.555 60.665 134.815 60.925 ;
        RECT 136.835 60.985 137.095 61.245 ;
        RECT 136.835 60.665 137.095 60.925 ;
        RECT 139.115 60.985 139.375 61.245 ;
        RECT 139.115 60.665 139.375 60.925 ;
        RECT 141.395 60.985 141.655 61.245 ;
        RECT 141.395 60.665 141.655 60.925 ;
        RECT 143.675 60.985 143.935 61.245 ;
        RECT 143.675 60.665 143.935 60.925 ;
        RECT 144.345 60.985 144.605 61.245 ;
        RECT 144.345 60.665 144.605 60.925 ;
        RECT 38.315 59.245 38.575 59.505 ;
        RECT 79.205 52.865 79.465 53.125 ;
        RECT 79.525 52.865 79.785 53.125 ;
        RECT 79.845 52.865 80.105 53.125 ;
        RECT 55.935 52.330 56.195 52.590 ;
        RECT 55.935 52.010 56.195 52.270 ;
        RECT 55.935 51.690 56.195 51.950 ;
        RECT 65.845 52.330 66.105 52.590 ;
        RECT 65.845 52.010 66.105 52.270 ;
        RECT 65.845 51.690 66.105 51.950 ;
        RECT 68.125 52.330 68.385 52.590 ;
        RECT 68.125 52.010 68.385 52.270 ;
        RECT 68.125 51.690 68.385 51.950 ;
        RECT 70.405 52.330 70.665 52.590 ;
        RECT 70.405 52.010 70.665 52.270 ;
        RECT 70.405 51.690 70.665 51.950 ;
        RECT 72.685 52.330 72.945 52.590 ;
        RECT 72.685 52.010 72.945 52.270 ;
        RECT 72.685 51.690 72.945 51.950 ;
        RECT 74.965 52.330 75.225 52.590 ;
        RECT 74.965 52.010 75.225 52.270 ;
        RECT 74.965 51.690 75.225 51.950 ;
        RECT 77.245 52.330 77.505 52.590 ;
        RECT 77.245 52.010 77.505 52.270 ;
        RECT 77.245 51.690 77.505 51.950 ;
        RECT 79.525 52.330 79.785 52.590 ;
        RECT 79.525 52.010 79.785 52.270 ;
        RECT 79.525 51.690 79.785 51.950 ;
        RECT 81.805 52.330 82.065 52.590 ;
        RECT 81.805 52.010 82.065 52.270 ;
        RECT 81.805 51.690 82.065 51.950 ;
        RECT 84.085 52.330 84.345 52.590 ;
        RECT 84.085 52.010 84.345 52.270 ;
        RECT 84.085 51.690 84.345 51.950 ;
        RECT 86.365 52.330 86.625 52.590 ;
        RECT 86.365 52.010 86.625 52.270 ;
        RECT 86.365 51.690 86.625 51.950 ;
        RECT 88.645 52.330 88.905 52.590 ;
        RECT 88.645 52.010 88.905 52.270 ;
        RECT 88.645 51.690 88.905 51.950 ;
        RECT 90.925 52.330 91.185 52.590 ;
        RECT 90.925 52.010 91.185 52.270 ;
        RECT 90.925 51.690 91.185 51.950 ;
        RECT 93.205 52.330 93.465 52.590 ;
        RECT 93.205 52.010 93.465 52.270 ;
        RECT 93.205 51.690 93.465 51.950 ;
        RECT 95.435 52.330 95.695 52.590 ;
        RECT 95.435 52.010 95.695 52.270 ;
        RECT 95.435 51.690 95.695 51.950 ;
        RECT 55.935 48.740 56.195 49.000 ;
        RECT 55.935 48.420 56.195 48.680 ;
        RECT 55.935 48.100 56.195 48.360 ;
        RECT 56.605 48.740 56.865 49.000 ;
        RECT 56.605 48.420 56.865 48.680 ;
        RECT 56.605 48.100 56.865 48.360 ;
        RECT 57.385 48.740 57.645 49.000 ;
        RECT 57.385 48.420 57.645 48.680 ;
        RECT 57.385 48.100 57.645 48.360 ;
        RECT 58.165 48.740 58.425 49.000 ;
        RECT 58.165 48.420 58.425 48.680 ;
        RECT 58.165 48.100 58.425 48.360 ;
        RECT 60.445 48.740 60.705 49.000 ;
        RECT 60.445 48.420 60.705 48.680 ;
        RECT 60.445 48.100 60.705 48.360 ;
        RECT 62.725 48.740 62.985 49.000 ;
        RECT 62.725 48.420 62.985 48.680 ;
        RECT 62.725 48.100 62.985 48.360 ;
        RECT 63.505 48.740 63.765 49.000 ;
        RECT 63.505 48.420 63.765 48.680 ;
        RECT 63.505 48.100 63.765 48.360 ;
        RECT 64.285 48.740 64.545 49.000 ;
        RECT 64.285 48.420 64.545 48.680 ;
        RECT 64.285 48.100 64.545 48.360 ;
        RECT 65.065 48.740 65.325 49.000 ;
        RECT 65.065 48.420 65.325 48.680 ;
        RECT 65.065 48.100 65.325 48.360 ;
        RECT 65.845 48.740 66.105 49.000 ;
        RECT 65.845 48.420 66.105 48.680 ;
        RECT 65.845 48.100 66.105 48.360 ;
        RECT 68.125 48.740 68.385 49.000 ;
        RECT 68.125 48.420 68.385 48.680 ;
        RECT 68.125 48.100 68.385 48.360 ;
        RECT 70.405 48.740 70.665 49.000 ;
        RECT 70.405 48.420 70.665 48.680 ;
        RECT 70.405 48.100 70.665 48.360 ;
        RECT 72.685 48.740 72.945 49.000 ;
        RECT 72.685 48.420 72.945 48.680 ;
        RECT 72.685 48.100 72.945 48.360 ;
        RECT 74.965 48.740 75.225 49.000 ;
        RECT 74.965 48.420 75.225 48.680 ;
        RECT 74.965 48.100 75.225 48.360 ;
        RECT 77.245 48.740 77.505 49.000 ;
        RECT 77.245 48.420 77.505 48.680 ;
        RECT 77.245 48.100 77.505 48.360 ;
        RECT 79.525 48.740 79.785 49.000 ;
        RECT 79.525 48.420 79.785 48.680 ;
        RECT 79.525 48.100 79.785 48.360 ;
        RECT 81.805 48.740 82.065 49.000 ;
        RECT 81.805 48.420 82.065 48.680 ;
        RECT 81.805 48.100 82.065 48.360 ;
        RECT 84.085 48.740 84.345 49.000 ;
        RECT 84.085 48.420 84.345 48.680 ;
        RECT 84.085 48.100 84.345 48.360 ;
        RECT 86.365 48.740 86.625 49.000 ;
        RECT 86.365 48.420 86.625 48.680 ;
        RECT 86.365 48.100 86.625 48.360 ;
        RECT 88.645 48.740 88.905 49.000 ;
        RECT 88.645 48.420 88.905 48.680 ;
        RECT 88.645 48.100 88.905 48.360 ;
        RECT 90.925 48.740 91.185 49.000 ;
        RECT 90.925 48.420 91.185 48.680 ;
        RECT 90.925 48.100 91.185 48.360 ;
        RECT 93.205 48.740 93.465 49.000 ;
        RECT 93.205 48.420 93.465 48.680 ;
        RECT 93.205 48.100 93.465 48.360 ;
        RECT 93.985 48.740 94.245 49.000 ;
        RECT 93.985 48.420 94.245 48.680 ;
        RECT 93.985 48.100 94.245 48.360 ;
        RECT 94.765 48.740 95.025 49.000 ;
        RECT 94.765 48.420 95.025 48.680 ;
        RECT 94.765 48.100 95.025 48.360 ;
        RECT 95.435 48.740 95.695 49.000 ;
        RECT 95.435 48.420 95.695 48.680 ;
        RECT 95.435 48.100 95.695 48.360 ;
        RECT 58.600 47.565 58.860 47.825 ;
        RECT 58.920 47.565 59.180 47.825 ;
        RECT 59.240 47.565 59.500 47.825 ;
        RECT 66.280 47.565 66.540 47.825 ;
        RECT 66.600 47.565 66.860 47.825 ;
        RECT 66.920 47.565 67.180 47.825 ;
        RECT 92.130 47.565 92.390 47.825 ;
        RECT 92.450 47.565 92.710 47.825 ;
        RECT 92.770 47.565 93.030 47.825 ;
        RECT 60.125 44.610 60.385 44.870 ;
        RECT 60.445 44.610 60.705 44.870 ;
        RECT 60.765 44.610 61.025 44.870 ;
        RECT 55.935 44.005 56.195 44.265 ;
        RECT 56.605 44.005 56.865 44.265 ;
        RECT 57.385 44.005 57.645 44.265 ;
        RECT 58.165 44.005 58.425 44.265 ;
        RECT 60.445 44.005 60.705 44.265 ;
        RECT 62.725 44.005 62.985 44.265 ;
        RECT 63.505 44.005 63.765 44.265 ;
        RECT 64.285 44.005 64.545 44.265 ;
        RECT 64.955 44.005 65.215 44.265 ;
        RECT 72.675 44.610 72.935 44.870 ;
        RECT 72.995 44.610 73.255 44.870 ;
        RECT 73.315 44.610 73.575 44.870 ;
        RECT 84.015 44.615 84.275 44.875 ;
        RECT 84.335 44.615 84.595 44.875 ;
        RECT 84.655 44.615 84.915 44.875 ;
        RECT 69.145 44.005 69.405 44.265 ;
        RECT 69.815 44.005 70.075 44.265 ;
        RECT 71.095 44.005 71.355 44.265 ;
        RECT 72.375 44.005 72.635 44.265 ;
        RECT 76.935 44.005 77.195 44.265 ;
        RECT 78.215 44.005 78.475 44.265 ;
        RECT 79.495 44.005 79.755 44.265 ;
        RECT 80.775 44.005 81.035 44.265 ;
        RECT 82.055 44.005 82.315 44.265 ;
        RECT 84.335 44.005 84.595 44.265 ;
        RECT 86.615 44.005 86.875 44.265 ;
        RECT 87.895 44.005 88.155 44.265 ;
        RECT 89.175 44.005 89.435 44.265 ;
        RECT 89.845 44.005 90.105 44.265 ;
        RECT 72.810 43.400 73.070 43.660 ;
        RECT 73.130 43.400 73.390 43.660 ;
        RECT 73.450 43.400 73.710 43.660 ;
        RECT 94.095 45.165 94.355 45.425 ;
        RECT 94.095 44.845 94.355 45.105 ;
        RECT 94.095 44.525 94.355 44.785 ;
        RECT 94.765 45.165 95.025 45.425 ;
        RECT 94.765 44.845 95.025 45.105 ;
        RECT 94.765 44.525 95.025 44.785 ;
        RECT 97.045 45.165 97.305 45.425 ;
        RECT 97.045 44.845 97.305 45.105 ;
        RECT 97.045 44.525 97.305 44.785 ;
        RECT 99.325 45.165 99.585 45.425 ;
        RECT 99.325 44.845 99.585 45.105 ;
        RECT 99.325 44.525 99.585 44.785 ;
        RECT 101.605 45.165 101.865 45.425 ;
        RECT 101.605 44.845 101.865 45.105 ;
        RECT 101.605 44.525 101.865 44.785 ;
        RECT 103.885 45.165 104.145 45.425 ;
        RECT 103.885 44.845 104.145 45.105 ;
        RECT 103.885 44.525 104.145 44.785 ;
        RECT 106.165 45.165 106.425 45.425 ;
        RECT 106.165 44.845 106.425 45.105 ;
        RECT 106.165 44.525 106.425 44.785 ;
        RECT 108.445 45.165 108.705 45.425 ;
        RECT 108.445 44.845 108.705 45.105 ;
        RECT 108.445 44.525 108.705 44.785 ;
        RECT 110.725 45.165 110.985 45.425 ;
        RECT 110.725 44.845 110.985 45.105 ;
        RECT 110.725 44.525 110.985 44.785 ;
        RECT 113.005 45.165 113.265 45.425 ;
        RECT 113.005 44.845 113.265 45.105 ;
        RECT 113.005 44.525 113.265 44.785 ;
        RECT 115.285 45.165 115.545 45.425 ;
        RECT 115.285 44.845 115.545 45.105 ;
        RECT 115.285 44.525 115.545 44.785 ;
        RECT 117.565 45.165 117.825 45.425 ;
        RECT 117.565 44.845 117.825 45.105 ;
        RECT 117.565 44.525 117.825 44.785 ;
        RECT 118.235 45.165 118.495 45.425 ;
        RECT 118.235 44.845 118.495 45.105 ;
        RECT 118.235 44.525 118.495 44.785 ;
        RECT 99.760 43.990 100.020 44.250 ;
        RECT 100.080 43.990 100.340 44.250 ;
        RECT 100.400 43.990 100.660 44.250 ;
        RECT 101.605 42.475 101.865 42.735 ;
        RECT 75.860 40.855 76.120 41.115 ;
        RECT 76.180 40.855 76.440 41.115 ;
        RECT 76.500 40.855 76.760 41.115 ;
        RECT 69.145 40.320 69.405 40.580 ;
        RECT 69.145 40.000 69.405 40.260 ;
        RECT 69.145 39.680 69.405 39.940 ;
        RECT 69.815 40.320 70.075 40.580 ;
        RECT 69.815 40.000 70.075 40.260 ;
        RECT 69.815 39.680 70.075 39.940 ;
        RECT 71.095 40.320 71.355 40.580 ;
        RECT 71.095 40.000 71.355 40.260 ;
        RECT 71.095 39.680 71.355 39.940 ;
        RECT 72.375 40.320 72.635 40.580 ;
        RECT 72.375 40.000 72.635 40.260 ;
        RECT 72.375 39.680 72.635 39.940 ;
        RECT 74.675 40.320 74.935 40.580 ;
        RECT 74.675 40.000 74.935 40.260 ;
        RECT 74.675 39.680 74.935 39.940 ;
        RECT 76.935 40.320 77.195 40.580 ;
        RECT 76.935 40.000 77.195 40.260 ;
        RECT 76.935 39.680 77.195 39.940 ;
        RECT 78.215 40.320 78.475 40.580 ;
        RECT 78.215 40.000 78.475 40.260 ;
        RECT 78.215 39.680 78.475 39.940 ;
        RECT 79.495 40.320 79.755 40.580 ;
        RECT 79.495 40.000 79.755 40.260 ;
        RECT 79.495 39.680 79.755 39.940 ;
        RECT 80.775 40.320 81.035 40.580 ;
        RECT 80.775 40.000 81.035 40.260 ;
        RECT 80.775 39.680 81.035 39.940 ;
        RECT 82.055 40.320 82.315 40.580 ;
        RECT 82.055 40.000 82.315 40.260 ;
        RECT 82.055 39.680 82.315 39.940 ;
        RECT 84.365 40.320 84.625 40.580 ;
        RECT 84.365 40.000 84.625 40.260 ;
        RECT 84.365 39.680 84.625 39.940 ;
        RECT 86.615 40.320 86.875 40.580 ;
        RECT 86.615 40.000 86.875 40.260 ;
        RECT 86.615 39.680 86.875 39.940 ;
        RECT 87.895 40.320 88.155 40.580 ;
        RECT 87.895 40.000 88.155 40.260 ;
        RECT 87.895 39.680 88.155 39.940 ;
        RECT 89.175 40.320 89.435 40.580 ;
        RECT 89.175 40.000 89.435 40.260 ;
        RECT 89.175 39.680 89.435 39.940 ;
        RECT 89.845 40.320 90.105 40.580 ;
        RECT 89.845 40.000 90.105 40.260 ;
        RECT 89.845 39.680 90.105 39.940 ;
        RECT 101.605 42.155 101.865 42.415 ;
        RECT 101.605 41.835 101.865 42.095 ;
        RECT 106.165 42.475 106.425 42.735 ;
        RECT 126.375 45.130 126.635 45.390 ;
        RECT 124.415 44.650 124.675 44.910 ;
        RECT 124.415 44.330 124.675 44.590 ;
        RECT 124.415 44.010 124.675 44.270 ;
        RECT 125.085 44.650 125.345 44.910 ;
        RECT 125.085 44.330 125.345 44.590 ;
        RECT 125.085 44.010 125.345 44.270 ;
        RECT 125.515 44.650 125.775 44.910 ;
        RECT 125.515 44.330 125.775 44.590 ;
        RECT 125.515 44.010 125.775 44.270 ;
        RECT 125.945 44.650 126.205 44.910 ;
        RECT 125.945 44.330 126.205 44.590 ;
        RECT 125.945 44.010 126.205 44.270 ;
        RECT 126.375 44.810 126.635 45.070 ;
        RECT 127.235 45.130 127.495 45.390 ;
        RECT 126.375 44.490 126.635 44.750 ;
        RECT 126.375 44.170 126.635 44.430 ;
        RECT 126.375 43.850 126.635 44.110 ;
        RECT 126.805 44.650 127.065 44.910 ;
        RECT 126.805 44.330 127.065 44.590 ;
        RECT 126.805 44.010 127.065 44.270 ;
        RECT 127.235 44.810 127.495 45.070 ;
        RECT 127.235 44.490 127.495 44.750 ;
        RECT 127.235 44.170 127.495 44.430 ;
        RECT 126.375 43.530 126.635 43.790 ;
        RECT 127.235 43.850 127.495 44.110 ;
        RECT 127.665 44.650 127.925 44.910 ;
        RECT 127.665 44.330 127.925 44.590 ;
        RECT 127.665 44.010 127.925 44.270 ;
        RECT 128.095 44.650 128.355 44.910 ;
        RECT 128.095 44.330 128.355 44.590 ;
        RECT 128.095 44.010 128.355 44.270 ;
        RECT 128.525 44.650 128.785 44.910 ;
        RECT 128.525 44.330 128.785 44.590 ;
        RECT 128.525 44.010 128.785 44.270 ;
        RECT 129.195 44.650 129.455 44.910 ;
        RECT 129.195 44.330 129.455 44.590 ;
        RECT 129.195 44.010 129.455 44.270 ;
        RECT 127.235 43.530 127.495 43.790 ;
        RECT 106.165 42.155 106.425 42.415 ;
        RECT 137.035 45.130 137.295 45.390 ;
        RECT 135.075 44.650 135.335 44.910 ;
        RECT 135.075 44.330 135.335 44.590 ;
        RECT 135.075 44.010 135.335 44.270 ;
        RECT 135.745 44.650 136.005 44.910 ;
        RECT 135.745 44.330 136.005 44.590 ;
        RECT 135.745 44.010 136.005 44.270 ;
        RECT 136.175 44.650 136.435 44.910 ;
        RECT 136.175 44.330 136.435 44.590 ;
        RECT 136.175 44.010 136.435 44.270 ;
        RECT 136.605 44.650 136.865 44.910 ;
        RECT 136.605 44.330 136.865 44.590 ;
        RECT 136.605 44.010 136.865 44.270 ;
        RECT 137.035 44.810 137.295 45.070 ;
        RECT 137.895 45.130 138.155 45.390 ;
        RECT 137.035 44.490 137.295 44.750 ;
        RECT 137.035 44.170 137.295 44.430 ;
        RECT 137.035 43.850 137.295 44.110 ;
        RECT 137.465 44.650 137.725 44.910 ;
        RECT 137.465 44.330 137.725 44.590 ;
        RECT 137.465 44.010 137.725 44.270 ;
        RECT 137.895 44.810 138.155 45.070 ;
        RECT 138.755 45.130 139.015 45.390 ;
        RECT 137.895 44.490 138.155 44.750 ;
        RECT 137.895 44.170 138.155 44.430 ;
        RECT 137.035 43.530 137.295 43.790 ;
        RECT 137.895 43.850 138.155 44.110 ;
        RECT 138.325 44.650 138.585 44.910 ;
        RECT 138.325 44.330 138.585 44.590 ;
        RECT 138.325 44.010 138.585 44.270 ;
        RECT 138.755 44.810 139.015 45.070 ;
        RECT 139.615 45.130 139.875 45.390 ;
        RECT 138.755 44.490 139.015 44.750 ;
        RECT 138.755 44.170 139.015 44.430 ;
        RECT 137.895 43.530 138.155 43.790 ;
        RECT 138.755 43.850 139.015 44.110 ;
        RECT 139.185 44.650 139.445 44.910 ;
        RECT 139.185 44.330 139.445 44.590 ;
        RECT 139.185 44.010 139.445 44.270 ;
        RECT 139.615 44.810 139.875 45.070 ;
        RECT 140.475 45.130 140.735 45.390 ;
        RECT 139.615 44.490 139.875 44.750 ;
        RECT 139.615 44.170 139.875 44.430 ;
        RECT 138.755 43.530 139.015 43.790 ;
        RECT 139.615 43.850 139.875 44.110 ;
        RECT 140.045 44.650 140.305 44.910 ;
        RECT 140.045 44.330 140.305 44.590 ;
        RECT 140.045 44.010 140.305 44.270 ;
        RECT 140.475 44.810 140.735 45.070 ;
        RECT 141.335 45.130 141.595 45.390 ;
        RECT 140.475 44.490 140.735 44.750 ;
        RECT 140.475 44.170 140.735 44.430 ;
        RECT 139.615 43.530 139.875 43.790 ;
        RECT 140.475 43.850 140.735 44.110 ;
        RECT 140.905 44.650 141.165 44.910 ;
        RECT 140.905 44.330 141.165 44.590 ;
        RECT 140.905 44.010 141.165 44.270 ;
        RECT 141.335 44.810 141.595 45.070 ;
        RECT 142.195 45.130 142.455 45.390 ;
        RECT 141.335 44.490 141.595 44.750 ;
        RECT 141.335 44.170 141.595 44.430 ;
        RECT 140.475 43.530 140.735 43.790 ;
        RECT 141.335 43.850 141.595 44.110 ;
        RECT 141.765 44.650 142.025 44.910 ;
        RECT 141.765 44.330 142.025 44.590 ;
        RECT 141.765 44.010 142.025 44.270 ;
        RECT 142.195 44.810 142.455 45.070 ;
        RECT 142.195 44.490 142.455 44.750 ;
        RECT 142.195 44.170 142.455 44.430 ;
        RECT 141.335 43.530 141.595 43.790 ;
        RECT 142.195 43.850 142.455 44.110 ;
        RECT 142.625 44.650 142.885 44.910 ;
        RECT 142.625 44.330 142.885 44.590 ;
        RECT 142.625 44.010 142.885 44.270 ;
        RECT 143.055 44.650 143.315 44.910 ;
        RECT 143.055 44.330 143.315 44.590 ;
        RECT 143.055 44.010 143.315 44.270 ;
        RECT 143.485 44.650 143.745 44.910 ;
        RECT 143.485 44.330 143.745 44.590 ;
        RECT 143.485 44.010 143.745 44.270 ;
        RECT 144.155 44.650 144.415 44.910 ;
        RECT 144.155 44.330 144.415 44.590 ;
        RECT 144.155 44.010 144.415 44.270 ;
        RECT 142.195 43.530 142.455 43.790 ;
        RECT 106.165 41.835 106.425 42.095 ;
        RECT 99.760 40.900 100.020 41.160 ;
        RECT 100.080 40.900 100.340 41.160 ;
        RECT 100.400 40.900 100.660 41.160 ;
        RECT 125.180 42.155 125.440 42.415 ;
        RECT 125.500 42.155 125.760 42.415 ;
        RECT 94.095 40.295 94.355 40.555 ;
        RECT 94.765 40.295 95.025 40.555 ;
        RECT 97.045 40.295 97.305 40.555 ;
        RECT 99.325 40.295 99.585 40.555 ;
        RECT 101.605 40.295 101.865 40.555 ;
        RECT 103.885 40.295 104.145 40.555 ;
        RECT 106.165 40.295 106.425 40.555 ;
        RECT 108.445 40.295 108.705 40.555 ;
        RECT 110.725 40.295 110.985 40.555 ;
        RECT 113.005 40.295 113.265 40.555 ;
        RECT 115.285 40.295 115.545 40.555 ;
        RECT 117.565 40.295 117.825 40.555 ;
        RECT 118.235 40.295 118.495 40.555 ;
        RECT 135.840 42.155 136.100 42.415 ;
        RECT 136.160 42.155 136.420 42.415 ;
        RECT 124.415 40.800 124.675 41.060 ;
        RECT 124.415 40.480 124.675 40.740 ;
        RECT 124.415 40.160 124.675 40.420 ;
        RECT 125.085 40.800 125.345 41.060 ;
        RECT 125.085 40.480 125.345 40.740 ;
        RECT 125.085 40.160 125.345 40.420 ;
        RECT 125.515 40.800 125.775 41.060 ;
        RECT 125.515 40.480 125.775 40.740 ;
        RECT 125.515 40.160 125.775 40.420 ;
        RECT 125.945 40.800 126.205 41.060 ;
        RECT 125.945 40.480 126.205 40.740 ;
        RECT 125.945 40.160 126.205 40.420 ;
        RECT 126.375 40.800 126.635 41.060 ;
        RECT 126.375 40.480 126.635 40.740 ;
        RECT 126.375 40.160 126.635 40.420 ;
        RECT 126.805 40.800 127.065 41.060 ;
        RECT 126.805 40.480 127.065 40.740 ;
        RECT 126.805 40.160 127.065 40.420 ;
        RECT 127.235 40.800 127.495 41.060 ;
        RECT 127.235 40.480 127.495 40.740 ;
        RECT 127.235 40.160 127.495 40.420 ;
        RECT 127.665 40.800 127.925 41.060 ;
        RECT 127.665 40.480 127.925 40.740 ;
        RECT 127.665 40.160 127.925 40.420 ;
        RECT 128.095 40.800 128.355 41.060 ;
        RECT 128.095 40.480 128.355 40.740 ;
        RECT 128.095 40.160 128.355 40.420 ;
        RECT 128.525 40.800 128.785 41.060 ;
        RECT 128.525 40.480 128.785 40.740 ;
        RECT 128.525 40.160 128.785 40.420 ;
        RECT 129.195 40.800 129.455 41.060 ;
        RECT 129.195 40.480 129.455 40.740 ;
        RECT 129.195 40.160 129.455 40.420 ;
        RECT 137.895 42.475 138.155 42.735 ;
        RECT 137.895 42.155 138.155 42.415 ;
        RECT 137.895 41.835 138.155 42.095 ;
        RECT 135.075 40.800 135.335 41.060 ;
        RECT 135.075 40.480 135.335 40.740 ;
        RECT 135.075 40.160 135.335 40.420 ;
        RECT 135.745 40.800 136.005 41.060 ;
        RECT 135.745 40.480 136.005 40.740 ;
        RECT 135.745 40.160 136.005 40.420 ;
        RECT 136.175 40.800 136.435 41.060 ;
        RECT 136.175 40.480 136.435 40.740 ;
        RECT 136.175 40.160 136.435 40.420 ;
        RECT 136.605 40.800 136.865 41.060 ;
        RECT 136.605 40.480 136.865 40.740 ;
        RECT 136.605 40.160 136.865 40.420 ;
        RECT 137.035 40.800 137.295 41.060 ;
        RECT 137.035 40.480 137.295 40.740 ;
        RECT 137.035 40.160 137.295 40.420 ;
        RECT 137.465 40.800 137.725 41.060 ;
        RECT 137.465 40.480 137.725 40.740 ;
        RECT 137.465 40.160 137.725 40.420 ;
        RECT 137.895 40.800 138.155 41.060 ;
        RECT 137.895 40.480 138.155 40.740 ;
        RECT 137.895 40.160 138.155 40.420 ;
        RECT 138.325 40.800 138.585 41.060 ;
        RECT 138.325 40.480 138.585 40.740 ;
        RECT 138.325 40.160 138.585 40.420 ;
        RECT 138.755 40.800 139.015 41.060 ;
        RECT 138.755 40.480 139.015 40.740 ;
        RECT 138.755 40.160 139.015 40.420 ;
        RECT 139.185 40.800 139.445 41.060 ;
        RECT 139.185 40.480 139.445 40.740 ;
        RECT 139.185 40.160 139.445 40.420 ;
        RECT 139.615 40.800 139.875 41.060 ;
        RECT 139.615 40.480 139.875 40.740 ;
        RECT 139.615 40.160 139.875 40.420 ;
        RECT 140.045 40.800 140.305 41.060 ;
        RECT 140.045 40.480 140.305 40.740 ;
        RECT 140.045 40.160 140.305 40.420 ;
        RECT 140.475 40.800 140.735 41.060 ;
        RECT 140.475 40.480 140.735 40.740 ;
        RECT 140.475 40.160 140.735 40.420 ;
        RECT 140.905 40.800 141.165 41.060 ;
        RECT 140.905 40.480 141.165 40.740 ;
        RECT 140.905 40.160 141.165 40.420 ;
        RECT 141.335 40.800 141.595 41.060 ;
        RECT 141.335 40.480 141.595 40.740 ;
        RECT 141.335 40.160 141.595 40.420 ;
        RECT 141.765 40.800 142.025 41.060 ;
        RECT 141.765 40.480 142.025 40.740 ;
        RECT 141.765 40.160 142.025 40.420 ;
        RECT 142.195 40.800 142.455 41.060 ;
        RECT 142.195 40.480 142.455 40.740 ;
        RECT 142.195 40.160 142.455 40.420 ;
        RECT 142.625 40.800 142.885 41.060 ;
        RECT 142.625 40.480 142.885 40.740 ;
        RECT 142.625 40.160 142.885 40.420 ;
        RECT 143.055 40.800 143.315 41.060 ;
        RECT 143.055 40.480 143.315 40.740 ;
        RECT 143.055 40.160 143.315 40.420 ;
        RECT 143.485 40.800 143.745 41.060 ;
        RECT 143.485 40.480 143.745 40.740 ;
        RECT 143.485 40.160 143.745 40.420 ;
        RECT 144.155 40.800 144.415 41.060 ;
        RECT 144.155 40.480 144.415 40.740 ;
        RECT 144.155 40.160 144.415 40.420 ;
        RECT 66.280 36.455 66.540 36.715 ;
        RECT 66.600 36.455 66.860 36.715 ;
        RECT 92.450 36.455 92.710 36.715 ;
        RECT 92.770 36.455 93.030 36.715 ;
        RECT 64.655 35.850 64.915 36.110 ;
        RECT 65.285 35.850 65.545 36.110 ;
        RECT 67.845 35.850 68.105 36.110 ;
        RECT 70.125 35.850 70.385 36.110 ;
        RECT 72.405 35.850 72.665 36.110 ;
        RECT 74.685 35.850 74.945 36.110 ;
        RECT 76.965 35.850 77.225 36.110 ;
        RECT 78.245 35.850 78.505 36.110 ;
        RECT 79.525 35.850 79.785 36.110 ;
        RECT 80.805 35.850 81.065 36.110 ;
        RECT 82.085 35.850 82.345 36.110 ;
        RECT 84.365 35.850 84.625 36.110 ;
        RECT 86.645 35.850 86.905 36.110 ;
        RECT 88.925 35.850 89.185 36.110 ;
        RECT 91.205 35.850 91.465 36.110 ;
        RECT 93.765 35.850 94.025 36.110 ;
        RECT 94.395 35.850 94.655 36.110 ;
        RECT 126.565 37.340 126.825 37.600 ;
        RECT 126.885 37.340 127.145 37.600 ;
        RECT 124.765 36.570 125.025 36.830 ;
        RECT 124.765 36.250 125.025 36.510 ;
        RECT 125.435 36.570 125.695 36.830 ;
        RECT 125.435 36.250 125.695 36.510 ;
        RECT 125.865 36.570 126.125 36.830 ;
        RECT 125.865 36.250 126.125 36.510 ;
        RECT 126.295 36.570 126.555 36.830 ;
        RECT 126.295 36.250 126.555 36.510 ;
        RECT 126.725 36.805 126.985 37.065 ;
        RECT 126.725 36.485 126.985 36.745 ;
        RECT 126.725 36.165 126.985 36.425 ;
        RECT 127.155 36.570 127.415 36.830 ;
        RECT 127.155 36.250 127.415 36.510 ;
        RECT 127.585 36.805 127.845 37.065 ;
        RECT 127.585 36.485 127.845 36.745 ;
        RECT 127.585 36.165 127.845 36.425 ;
        RECT 128.015 36.570 128.275 36.830 ;
        RECT 128.015 36.250 128.275 36.510 ;
        RECT 128.445 36.570 128.705 36.830 ;
        RECT 128.445 36.250 128.705 36.510 ;
        RECT 128.875 36.570 129.135 36.830 ;
        RECT 128.875 36.250 129.135 36.510 ;
        RECT 129.525 36.570 129.785 36.830 ;
        RECT 129.525 36.250 129.785 36.510 ;
        RECT 135.075 36.830 135.335 37.090 ;
        RECT 135.075 36.510 135.335 36.770 ;
        RECT 135.075 36.190 135.335 36.450 ;
        RECT 135.745 36.830 136.005 37.090 ;
        RECT 135.745 36.510 136.005 36.770 ;
        RECT 135.745 36.190 136.005 36.450 ;
        RECT 136.175 36.830 136.435 37.090 ;
        RECT 136.175 36.510 136.435 36.770 ;
        RECT 136.175 36.190 136.435 36.450 ;
        RECT 136.605 36.830 136.865 37.090 ;
        RECT 136.605 36.510 136.865 36.770 ;
        RECT 136.605 36.190 136.865 36.450 ;
        RECT 137.035 36.830 137.295 37.090 ;
        RECT 137.035 36.510 137.295 36.770 ;
        RECT 137.035 36.190 137.295 36.450 ;
        RECT 137.465 36.830 137.725 37.090 ;
        RECT 137.465 36.510 137.725 36.770 ;
        RECT 137.465 36.190 137.725 36.450 ;
        RECT 137.895 36.830 138.155 37.090 ;
        RECT 137.895 36.510 138.155 36.770 ;
        RECT 137.895 36.190 138.155 36.450 ;
        RECT 138.325 36.830 138.585 37.090 ;
        RECT 138.325 36.510 138.585 36.770 ;
        RECT 138.325 36.190 138.585 36.450 ;
        RECT 138.755 36.830 139.015 37.090 ;
        RECT 138.755 36.510 139.015 36.770 ;
        RECT 138.755 36.190 139.015 36.450 ;
        RECT 139.185 36.830 139.445 37.090 ;
        RECT 139.185 36.510 139.445 36.770 ;
        RECT 139.185 36.190 139.445 36.450 ;
        RECT 139.615 36.830 139.875 37.090 ;
        RECT 139.615 36.510 139.875 36.770 ;
        RECT 139.615 36.190 139.875 36.450 ;
        RECT 140.045 36.830 140.305 37.090 ;
        RECT 140.045 36.510 140.305 36.770 ;
        RECT 140.045 36.190 140.305 36.450 ;
        RECT 140.475 36.830 140.735 37.090 ;
        RECT 140.475 36.510 140.735 36.770 ;
        RECT 140.475 36.190 140.735 36.450 ;
        RECT 140.905 36.830 141.165 37.090 ;
        RECT 140.905 36.510 141.165 36.770 ;
        RECT 140.905 36.190 141.165 36.450 ;
        RECT 141.335 36.830 141.595 37.090 ;
        RECT 141.335 36.510 141.595 36.770 ;
        RECT 141.335 36.190 141.595 36.450 ;
        RECT 141.765 36.830 142.025 37.090 ;
        RECT 141.765 36.510 142.025 36.770 ;
        RECT 141.765 36.190 142.025 36.450 ;
        RECT 142.195 36.830 142.455 37.090 ;
        RECT 142.195 36.510 142.455 36.770 ;
        RECT 142.195 36.190 142.455 36.450 ;
        RECT 142.625 36.830 142.885 37.090 ;
        RECT 142.625 36.510 142.885 36.770 ;
        RECT 142.625 36.190 142.885 36.450 ;
        RECT 143.055 36.830 143.315 37.090 ;
        RECT 143.055 36.510 143.315 36.770 ;
        RECT 143.055 36.190 143.315 36.450 ;
        RECT 143.485 36.830 143.745 37.090 ;
        RECT 143.485 36.510 143.745 36.770 ;
        RECT 143.485 36.190 143.745 36.450 ;
        RECT 144.155 36.830 144.415 37.090 ;
        RECT 144.155 36.510 144.415 36.770 ;
        RECT 144.155 36.190 144.415 36.450 ;
        RECT 125.645 34.835 125.905 35.095 ;
        RECT 125.965 34.835 126.225 35.095 ;
        RECT 135.840 34.835 136.100 35.095 ;
        RECT 136.160 34.835 136.420 35.095 ;
        RECT 64.655 33.110 64.915 33.370 ;
        RECT 65.685 33.110 65.945 33.370 ;
        RECT 68.965 33.110 69.225 33.370 ;
        RECT 72.245 33.110 72.505 33.370 ;
        RECT 79.525 33.110 79.785 33.370 ;
        RECT 86.805 33.110 87.065 33.370 ;
        RECT 90.085 33.110 90.345 33.370 ;
        RECT 93.365 33.110 93.625 33.370 ;
        RECT 94.395 33.110 94.655 33.370 ;
        RECT 80.605 32.505 80.865 32.765 ;
        RECT 80.925 32.505 81.185 32.765 ;
        RECT 81.245 32.505 81.505 32.765 ;
        RECT 81.565 32.505 81.825 32.765 ;
        RECT 124.765 33.345 125.025 33.605 ;
        RECT 124.765 33.025 125.025 33.285 ;
        RECT 125.435 33.345 125.695 33.605 ;
        RECT 125.435 33.025 125.695 33.285 ;
        RECT 125.865 33.345 126.125 33.605 ;
        RECT 125.865 33.025 126.125 33.285 ;
        RECT 126.295 33.505 126.555 33.765 ;
        RECT 126.295 33.185 126.555 33.445 ;
        RECT 126.295 32.865 126.555 33.125 ;
        RECT 126.725 33.505 126.985 33.765 ;
        RECT 126.725 33.185 126.985 33.445 ;
        RECT 126.725 32.865 126.985 33.125 ;
        RECT 127.155 33.505 127.415 33.765 ;
        RECT 127.155 33.185 127.415 33.445 ;
        RECT 127.155 32.865 127.415 33.125 ;
        RECT 127.585 33.505 127.845 33.765 ;
        RECT 127.585 33.185 127.845 33.445 ;
        RECT 127.585 32.865 127.845 33.125 ;
        RECT 128.015 33.505 128.275 33.765 ;
        RECT 128.015 33.185 128.275 33.445 ;
        RECT 128.015 32.865 128.275 33.125 ;
        RECT 128.445 33.345 128.705 33.605 ;
        RECT 128.445 33.025 128.705 33.285 ;
        RECT 128.875 33.345 129.135 33.605 ;
        RECT 128.875 33.025 129.135 33.285 ;
        RECT 129.525 33.345 129.785 33.605 ;
        RECT 129.525 33.025 129.785 33.285 ;
        RECT 124.765 31.770 125.025 32.030 ;
        RECT 124.765 31.450 125.025 31.710 ;
        RECT 125.435 31.770 125.695 32.030 ;
        RECT 125.435 31.450 125.695 31.710 ;
        RECT 125.865 31.770 126.125 32.030 ;
        RECT 125.865 31.450 126.125 31.710 ;
        RECT 126.295 31.770 126.555 32.030 ;
        RECT 126.295 31.450 126.555 31.710 ;
        RECT 126.725 31.855 126.985 32.115 ;
        RECT 126.725 31.535 126.985 31.795 ;
        RECT 126.725 31.215 126.985 31.475 ;
        RECT 127.155 31.770 127.415 32.030 ;
        RECT 127.155 31.450 127.415 31.710 ;
        RECT 127.585 31.855 127.845 32.115 ;
        RECT 127.585 31.535 127.845 31.795 ;
        RECT 127.585 31.215 127.845 31.475 ;
        RECT 128.015 31.770 128.275 32.030 ;
        RECT 128.015 31.450 128.275 31.710 ;
        RECT 128.445 31.770 128.705 32.030 ;
        RECT 128.445 31.450 128.705 31.710 ;
        RECT 128.875 31.770 129.135 32.030 ;
        RECT 128.875 31.450 129.135 31.710 ;
        RECT 129.525 31.770 129.785 32.030 ;
        RECT 129.525 31.450 129.785 31.710 ;
        RECT 126.675 30.680 126.935 30.940 ;
        RECT 126.995 30.680 127.255 30.940 ;
        RECT 127.315 30.680 127.575 30.940 ;
        RECT 127.635 30.680 127.895 30.940 ;
        RECT 126.675 29.620 126.935 29.880 ;
        RECT 126.995 29.620 127.255 29.880 ;
        RECT 127.315 29.620 127.575 29.880 ;
        RECT 127.635 29.620 127.895 29.880 ;
        RECT 124.765 28.850 125.025 29.110 ;
        RECT 80.605 28.025 80.865 28.285 ;
        RECT 80.925 28.025 81.185 28.285 ;
        RECT 81.245 28.025 81.505 28.285 ;
        RECT 81.565 28.025 81.825 28.285 ;
        RECT 64.655 27.420 64.915 27.680 ;
        RECT 65.685 27.420 65.945 27.680 ;
        RECT 68.965 27.420 69.225 27.680 ;
        RECT 72.245 27.420 72.505 27.680 ;
        RECT 79.525 27.420 79.785 27.680 ;
        RECT 86.805 27.420 87.065 27.680 ;
        RECT 90.085 27.420 90.345 27.680 ;
        RECT 93.365 27.420 93.625 27.680 ;
        RECT 94.395 27.420 94.655 27.680 ;
        RECT 124.765 28.530 125.025 28.790 ;
        RECT 125.435 28.850 125.695 29.110 ;
        RECT 125.435 28.530 125.695 28.790 ;
        RECT 125.865 28.850 126.125 29.110 ;
        RECT 125.865 28.530 126.125 28.790 ;
        RECT 126.295 28.850 126.555 29.110 ;
        RECT 126.295 28.530 126.555 28.790 ;
        RECT 126.725 29.085 126.985 29.345 ;
        RECT 126.725 28.765 126.985 29.025 ;
        RECT 126.725 28.445 126.985 28.705 ;
        RECT 127.155 28.850 127.415 29.110 ;
        RECT 127.155 28.530 127.415 28.790 ;
        RECT 127.585 29.085 127.845 29.345 ;
        RECT 127.585 28.765 127.845 29.025 ;
        RECT 127.585 28.445 127.845 28.705 ;
        RECT 128.015 28.850 128.275 29.110 ;
        RECT 128.015 28.530 128.275 28.790 ;
        RECT 128.445 28.850 128.705 29.110 ;
        RECT 128.445 28.530 128.705 28.790 ;
        RECT 128.875 28.850 129.135 29.110 ;
        RECT 128.875 28.530 129.135 28.790 ;
        RECT 129.525 28.850 129.785 29.110 ;
        RECT 129.525 28.530 129.785 28.790 ;
        RECT 124.765 27.275 125.025 27.535 ;
        RECT 124.765 26.955 125.025 27.215 ;
        RECT 125.435 27.275 125.695 27.535 ;
        RECT 125.435 26.955 125.695 27.215 ;
        RECT 125.865 27.275 126.125 27.535 ;
        RECT 125.865 26.955 126.125 27.215 ;
        RECT 126.295 27.435 126.555 27.695 ;
        RECT 126.295 27.115 126.555 27.375 ;
        RECT 126.295 26.795 126.555 27.055 ;
        RECT 126.725 27.435 126.985 27.695 ;
        RECT 126.725 27.115 126.985 27.375 ;
        RECT 126.725 26.795 126.985 27.055 ;
        RECT 127.155 27.435 127.415 27.695 ;
        RECT 127.155 27.115 127.415 27.375 ;
        RECT 127.155 26.795 127.415 27.055 ;
        RECT 127.585 27.435 127.845 27.695 ;
        RECT 127.585 27.115 127.845 27.375 ;
        RECT 127.585 26.795 127.845 27.055 ;
        RECT 128.015 27.435 128.275 27.695 ;
        RECT 137.895 35.155 138.155 35.415 ;
        RECT 137.895 34.835 138.155 35.095 ;
        RECT 137.895 34.515 138.155 34.775 ;
        RECT 137.035 33.460 137.295 33.720 ;
        RECT 135.075 32.980 135.335 33.240 ;
        RECT 135.075 32.660 135.335 32.920 ;
        RECT 135.075 32.340 135.335 32.600 ;
        RECT 135.745 32.980 136.005 33.240 ;
        RECT 135.745 32.660 136.005 32.920 ;
        RECT 135.745 32.340 136.005 32.600 ;
        RECT 136.175 32.980 136.435 33.240 ;
        RECT 136.175 32.660 136.435 32.920 ;
        RECT 136.175 32.340 136.435 32.600 ;
        RECT 136.605 32.980 136.865 33.240 ;
        RECT 136.605 32.660 136.865 32.920 ;
        RECT 136.605 32.340 136.865 32.600 ;
        RECT 137.035 33.140 137.295 33.400 ;
        RECT 137.895 33.460 138.155 33.720 ;
        RECT 137.035 32.820 137.295 33.080 ;
        RECT 137.035 32.500 137.295 32.760 ;
        RECT 137.035 32.180 137.295 32.440 ;
        RECT 137.465 32.980 137.725 33.240 ;
        RECT 137.465 32.660 137.725 32.920 ;
        RECT 137.465 32.340 137.725 32.600 ;
        RECT 137.895 33.140 138.155 33.400 ;
        RECT 138.755 33.460 139.015 33.720 ;
        RECT 137.895 32.820 138.155 33.080 ;
        RECT 137.895 32.500 138.155 32.760 ;
        RECT 137.035 31.860 137.295 32.120 ;
        RECT 137.895 32.180 138.155 32.440 ;
        RECT 138.325 32.980 138.585 33.240 ;
        RECT 138.325 32.660 138.585 32.920 ;
        RECT 138.325 32.340 138.585 32.600 ;
        RECT 138.755 33.140 139.015 33.400 ;
        RECT 139.615 33.460 139.875 33.720 ;
        RECT 138.755 32.820 139.015 33.080 ;
        RECT 138.755 32.500 139.015 32.760 ;
        RECT 137.895 31.860 138.155 32.120 ;
        RECT 138.755 32.180 139.015 32.440 ;
        RECT 139.185 32.980 139.445 33.240 ;
        RECT 139.185 32.660 139.445 32.920 ;
        RECT 139.185 32.340 139.445 32.600 ;
        RECT 139.615 33.140 139.875 33.400 ;
        RECT 140.475 33.460 140.735 33.720 ;
        RECT 139.615 32.820 139.875 33.080 ;
        RECT 139.615 32.500 139.875 32.760 ;
        RECT 138.755 31.860 139.015 32.120 ;
        RECT 139.615 32.180 139.875 32.440 ;
        RECT 140.045 32.980 140.305 33.240 ;
        RECT 140.045 32.660 140.305 32.920 ;
        RECT 140.045 32.340 140.305 32.600 ;
        RECT 140.475 33.140 140.735 33.400 ;
        RECT 141.335 33.460 141.595 33.720 ;
        RECT 140.475 32.820 140.735 33.080 ;
        RECT 140.475 32.500 140.735 32.760 ;
        RECT 139.615 31.860 139.875 32.120 ;
        RECT 140.475 32.180 140.735 32.440 ;
        RECT 140.905 32.980 141.165 33.240 ;
        RECT 140.905 32.660 141.165 32.920 ;
        RECT 140.905 32.340 141.165 32.600 ;
        RECT 141.335 33.140 141.595 33.400 ;
        RECT 142.195 33.460 142.455 33.720 ;
        RECT 141.335 32.820 141.595 33.080 ;
        RECT 141.335 32.500 141.595 32.760 ;
        RECT 140.475 31.860 140.735 32.120 ;
        RECT 141.335 32.180 141.595 32.440 ;
        RECT 141.765 32.980 142.025 33.240 ;
        RECT 141.765 32.660 142.025 32.920 ;
        RECT 141.765 32.340 142.025 32.600 ;
        RECT 142.195 33.140 142.455 33.400 ;
        RECT 142.195 32.820 142.455 33.080 ;
        RECT 142.195 32.500 142.455 32.760 ;
        RECT 141.335 31.860 141.595 32.120 ;
        RECT 142.195 32.180 142.455 32.440 ;
        RECT 142.625 32.980 142.885 33.240 ;
        RECT 142.625 32.660 142.885 32.920 ;
        RECT 142.625 32.340 142.885 32.600 ;
        RECT 143.055 32.980 143.315 33.240 ;
        RECT 143.055 32.660 143.315 32.920 ;
        RECT 143.055 32.340 143.315 32.600 ;
        RECT 143.485 32.980 143.745 33.240 ;
        RECT 143.485 32.660 143.745 32.920 ;
        RECT 143.485 32.340 143.745 32.600 ;
        RECT 144.155 32.980 144.415 33.240 ;
        RECT 144.155 32.660 144.415 32.920 ;
        RECT 144.155 32.340 144.415 32.600 ;
        RECT 142.195 31.860 142.455 32.120 ;
        RECT 137.035 30.370 137.295 30.630 ;
        RECT 135.075 29.890 135.335 30.150 ;
        RECT 135.075 29.570 135.335 29.830 ;
        RECT 135.075 29.250 135.335 29.510 ;
        RECT 135.745 29.890 136.005 30.150 ;
        RECT 135.745 29.570 136.005 29.830 ;
        RECT 135.745 29.250 136.005 29.510 ;
        RECT 136.175 29.890 136.435 30.150 ;
        RECT 136.175 29.570 136.435 29.830 ;
        RECT 136.175 29.250 136.435 29.510 ;
        RECT 136.605 29.890 136.865 30.150 ;
        RECT 136.605 29.570 136.865 29.830 ;
        RECT 136.605 29.250 136.865 29.510 ;
        RECT 137.035 30.050 137.295 30.310 ;
        RECT 137.895 30.370 138.155 30.630 ;
        RECT 137.035 29.730 137.295 29.990 ;
        RECT 137.035 29.410 137.295 29.670 ;
        RECT 137.035 29.090 137.295 29.350 ;
        RECT 137.465 29.890 137.725 30.150 ;
        RECT 137.465 29.570 137.725 29.830 ;
        RECT 137.465 29.250 137.725 29.510 ;
        RECT 137.895 30.050 138.155 30.310 ;
        RECT 138.755 30.370 139.015 30.630 ;
        RECT 137.895 29.730 138.155 29.990 ;
        RECT 137.895 29.410 138.155 29.670 ;
        RECT 137.035 28.770 137.295 29.030 ;
        RECT 137.895 29.090 138.155 29.350 ;
        RECT 138.325 29.890 138.585 30.150 ;
        RECT 138.325 29.570 138.585 29.830 ;
        RECT 138.325 29.250 138.585 29.510 ;
        RECT 138.755 30.050 139.015 30.310 ;
        RECT 139.615 30.370 139.875 30.630 ;
        RECT 138.755 29.730 139.015 29.990 ;
        RECT 138.755 29.410 139.015 29.670 ;
        RECT 137.895 28.770 138.155 29.030 ;
        RECT 138.755 29.090 139.015 29.350 ;
        RECT 139.185 29.890 139.445 30.150 ;
        RECT 139.185 29.570 139.445 29.830 ;
        RECT 139.185 29.250 139.445 29.510 ;
        RECT 139.615 30.050 139.875 30.310 ;
        RECT 140.475 30.370 140.735 30.630 ;
        RECT 139.615 29.730 139.875 29.990 ;
        RECT 139.615 29.410 139.875 29.670 ;
        RECT 138.755 28.770 139.015 29.030 ;
        RECT 139.615 29.090 139.875 29.350 ;
        RECT 140.045 29.890 140.305 30.150 ;
        RECT 140.045 29.570 140.305 29.830 ;
        RECT 140.045 29.250 140.305 29.510 ;
        RECT 140.475 30.050 140.735 30.310 ;
        RECT 141.335 30.370 141.595 30.630 ;
        RECT 140.475 29.730 140.735 29.990 ;
        RECT 140.475 29.410 140.735 29.670 ;
        RECT 139.615 28.770 139.875 29.030 ;
        RECT 140.475 29.090 140.735 29.350 ;
        RECT 140.905 29.890 141.165 30.150 ;
        RECT 140.905 29.570 141.165 29.830 ;
        RECT 140.905 29.250 141.165 29.510 ;
        RECT 141.335 30.050 141.595 30.310 ;
        RECT 142.195 30.370 142.455 30.630 ;
        RECT 141.335 29.730 141.595 29.990 ;
        RECT 141.335 29.410 141.595 29.670 ;
        RECT 140.475 28.770 140.735 29.030 ;
        RECT 141.335 29.090 141.595 29.350 ;
        RECT 141.765 29.890 142.025 30.150 ;
        RECT 141.765 29.570 142.025 29.830 ;
        RECT 141.765 29.250 142.025 29.510 ;
        RECT 142.195 30.050 142.455 30.310 ;
        RECT 142.195 29.730 142.455 29.990 ;
        RECT 142.195 29.410 142.455 29.670 ;
        RECT 141.335 28.770 141.595 29.030 ;
        RECT 142.195 29.090 142.455 29.350 ;
        RECT 142.625 29.890 142.885 30.150 ;
        RECT 142.625 29.570 142.885 29.830 ;
        RECT 142.625 29.250 142.885 29.510 ;
        RECT 143.055 29.890 143.315 30.150 ;
        RECT 143.055 29.570 143.315 29.830 ;
        RECT 143.055 29.250 143.315 29.510 ;
        RECT 143.485 29.890 143.745 30.150 ;
        RECT 143.485 29.570 143.745 29.830 ;
        RECT 143.485 29.250 143.745 29.510 ;
        RECT 144.155 29.890 144.415 30.150 ;
        RECT 144.155 29.570 144.415 29.830 ;
        RECT 144.155 29.250 144.415 29.510 ;
        RECT 142.195 28.770 142.455 29.030 ;
        RECT 128.015 27.115 128.275 27.375 ;
        RECT 128.015 26.795 128.275 27.055 ;
        RECT 128.445 27.275 128.705 27.535 ;
        RECT 128.445 26.955 128.705 27.215 ;
        RECT 128.875 27.275 129.135 27.535 ;
        RECT 128.875 26.955 129.135 27.215 ;
        RECT 129.525 27.275 129.785 27.535 ;
        RECT 135.840 27.395 136.100 27.655 ;
        RECT 136.160 27.395 136.420 27.655 ;
        RECT 129.525 26.955 129.785 27.215 ;
        RECT 137.895 27.715 138.155 27.975 ;
        RECT 137.895 27.395 138.155 27.655 ;
        RECT 137.895 27.075 138.155 27.335 ;
        RECT 135.075 26.040 135.335 26.300 ;
        RECT 125.645 25.465 125.905 25.725 ;
        RECT 125.965 25.465 126.225 25.725 ;
        RECT 64.655 24.680 64.915 24.940 ;
        RECT 65.285 24.680 65.545 24.940 ;
        RECT 67.845 24.680 68.105 24.940 ;
        RECT 70.125 24.680 70.385 24.940 ;
        RECT 72.405 24.680 72.665 24.940 ;
        RECT 74.685 24.680 74.945 24.940 ;
        RECT 76.965 24.680 77.225 24.940 ;
        RECT 78.245 24.680 78.505 24.940 ;
        RECT 79.525 24.680 79.785 24.940 ;
        RECT 80.805 24.680 81.065 24.940 ;
        RECT 82.085 24.680 82.345 24.940 ;
        RECT 84.365 24.680 84.625 24.940 ;
        RECT 86.645 24.680 86.905 24.940 ;
        RECT 88.925 24.680 89.185 24.940 ;
        RECT 91.205 24.680 91.465 24.940 ;
        RECT 93.765 24.680 94.025 24.940 ;
        RECT 94.395 24.680 94.655 24.940 ;
        RECT 66.280 24.075 66.540 24.335 ;
        RECT 66.600 24.075 66.860 24.335 ;
        RECT 92.450 24.075 92.710 24.335 ;
        RECT 92.770 24.075 93.030 24.335 ;
        RECT 135.075 25.720 135.335 25.980 ;
        RECT 135.075 25.400 135.335 25.660 ;
        RECT 135.745 26.040 136.005 26.300 ;
        RECT 135.745 25.720 136.005 25.980 ;
        RECT 135.745 25.400 136.005 25.660 ;
        RECT 136.175 26.040 136.435 26.300 ;
        RECT 136.175 25.720 136.435 25.980 ;
        RECT 136.175 25.400 136.435 25.660 ;
        RECT 136.605 26.040 136.865 26.300 ;
        RECT 136.605 25.720 136.865 25.980 ;
        RECT 136.605 25.400 136.865 25.660 ;
        RECT 137.035 26.040 137.295 26.300 ;
        RECT 137.035 25.720 137.295 25.980 ;
        RECT 137.035 25.400 137.295 25.660 ;
        RECT 137.465 26.040 137.725 26.300 ;
        RECT 137.465 25.720 137.725 25.980 ;
        RECT 137.465 25.400 137.725 25.660 ;
        RECT 137.895 26.040 138.155 26.300 ;
        RECT 137.895 25.720 138.155 25.980 ;
        RECT 137.895 25.400 138.155 25.660 ;
        RECT 138.325 26.040 138.585 26.300 ;
        RECT 138.325 25.720 138.585 25.980 ;
        RECT 138.325 25.400 138.585 25.660 ;
        RECT 138.755 26.040 139.015 26.300 ;
        RECT 138.755 25.720 139.015 25.980 ;
        RECT 138.755 25.400 139.015 25.660 ;
        RECT 139.185 26.040 139.445 26.300 ;
        RECT 139.185 25.720 139.445 25.980 ;
        RECT 139.185 25.400 139.445 25.660 ;
        RECT 139.615 26.040 139.875 26.300 ;
        RECT 139.615 25.720 139.875 25.980 ;
        RECT 139.615 25.400 139.875 25.660 ;
        RECT 140.045 26.040 140.305 26.300 ;
        RECT 140.045 25.720 140.305 25.980 ;
        RECT 140.045 25.400 140.305 25.660 ;
        RECT 140.475 26.040 140.735 26.300 ;
        RECT 140.475 25.720 140.735 25.980 ;
        RECT 140.475 25.400 140.735 25.660 ;
        RECT 140.905 26.040 141.165 26.300 ;
        RECT 140.905 25.720 141.165 25.980 ;
        RECT 140.905 25.400 141.165 25.660 ;
        RECT 141.335 26.040 141.595 26.300 ;
        RECT 141.335 25.720 141.595 25.980 ;
        RECT 141.335 25.400 141.595 25.660 ;
        RECT 141.765 26.040 142.025 26.300 ;
        RECT 141.765 25.720 142.025 25.980 ;
        RECT 141.765 25.400 142.025 25.660 ;
        RECT 142.195 26.040 142.455 26.300 ;
        RECT 142.195 25.720 142.455 25.980 ;
        RECT 142.195 25.400 142.455 25.660 ;
        RECT 142.625 26.040 142.885 26.300 ;
        RECT 142.625 25.720 142.885 25.980 ;
        RECT 142.625 25.400 142.885 25.660 ;
        RECT 143.055 26.040 143.315 26.300 ;
        RECT 143.055 25.720 143.315 25.980 ;
        RECT 143.055 25.400 143.315 25.660 ;
        RECT 143.485 26.040 143.745 26.300 ;
        RECT 143.485 25.720 143.745 25.980 ;
        RECT 143.485 25.400 143.745 25.660 ;
        RECT 144.155 26.040 144.415 26.300 ;
        RECT 144.155 25.720 144.415 25.980 ;
        RECT 144.155 25.400 144.415 25.660 ;
        RECT 124.765 24.050 125.025 24.310 ;
        RECT 124.765 23.730 125.025 23.990 ;
        RECT 125.435 24.050 125.695 24.310 ;
        RECT 125.435 23.730 125.695 23.990 ;
        RECT 125.865 24.050 126.125 24.310 ;
        RECT 125.865 23.730 126.125 23.990 ;
        RECT 126.295 24.050 126.555 24.310 ;
        RECT 126.295 23.730 126.555 23.990 ;
        RECT 126.725 24.135 126.985 24.395 ;
        RECT 126.725 23.815 126.985 24.075 ;
        RECT 126.725 23.495 126.985 23.755 ;
        RECT 127.155 24.050 127.415 24.310 ;
        RECT 127.155 23.730 127.415 23.990 ;
        RECT 127.585 24.135 127.845 24.395 ;
        RECT 127.585 23.815 127.845 24.075 ;
        RECT 127.585 23.495 127.845 23.755 ;
        RECT 128.015 24.050 128.275 24.310 ;
        RECT 128.015 23.730 128.275 23.990 ;
        RECT 128.445 24.050 128.705 24.310 ;
        RECT 128.445 23.730 128.705 23.990 ;
        RECT 128.875 24.050 129.135 24.310 ;
        RECT 128.875 23.730 129.135 23.990 ;
        RECT 129.525 24.050 129.785 24.310 ;
        RECT 129.525 23.730 129.785 23.990 ;
        RECT 126.565 22.960 126.825 23.220 ;
        RECT 126.885 22.960 127.145 23.220 ;
        RECT 69.145 20.850 69.405 21.110 ;
        RECT 69.145 20.530 69.405 20.790 ;
        RECT 69.145 20.210 69.405 20.470 ;
        RECT 69.815 20.850 70.075 21.110 ;
        RECT 69.815 20.530 70.075 20.790 ;
        RECT 69.815 20.210 70.075 20.470 ;
        RECT 71.095 20.850 71.355 21.110 ;
        RECT 71.095 20.530 71.355 20.790 ;
        RECT 71.095 20.210 71.355 20.470 ;
        RECT 72.375 20.850 72.635 21.110 ;
        RECT 72.375 20.530 72.635 20.790 ;
        RECT 72.375 20.210 72.635 20.470 ;
        RECT 74.675 20.850 74.935 21.110 ;
        RECT 74.675 20.530 74.935 20.790 ;
        RECT 74.675 20.210 74.935 20.470 ;
        RECT 76.935 20.850 77.195 21.110 ;
        RECT 76.935 20.530 77.195 20.790 ;
        RECT 76.935 20.210 77.195 20.470 ;
        RECT 78.215 20.850 78.475 21.110 ;
        RECT 78.215 20.530 78.475 20.790 ;
        RECT 78.215 20.210 78.475 20.470 ;
        RECT 79.495 20.850 79.755 21.110 ;
        RECT 79.495 20.530 79.755 20.790 ;
        RECT 79.495 20.210 79.755 20.470 ;
        RECT 80.775 20.850 81.035 21.110 ;
        RECT 80.775 20.530 81.035 20.790 ;
        RECT 80.775 20.210 81.035 20.470 ;
        RECT 82.055 20.850 82.315 21.110 ;
        RECT 82.055 20.530 82.315 20.790 ;
        RECT 82.055 20.210 82.315 20.470 ;
        RECT 84.365 20.850 84.625 21.110 ;
        RECT 84.365 20.530 84.625 20.790 ;
        RECT 84.365 20.210 84.625 20.470 ;
        RECT 86.615 20.850 86.875 21.110 ;
        RECT 86.615 20.530 86.875 20.790 ;
        RECT 86.615 20.210 86.875 20.470 ;
        RECT 87.895 20.850 88.155 21.110 ;
        RECT 87.895 20.530 88.155 20.790 ;
        RECT 87.895 20.210 88.155 20.470 ;
        RECT 89.175 20.850 89.435 21.110 ;
        RECT 89.175 20.530 89.435 20.790 ;
        RECT 89.175 20.210 89.435 20.470 ;
        RECT 89.845 20.850 90.105 21.110 ;
        RECT 89.845 20.530 90.105 20.790 ;
        RECT 89.845 20.210 90.105 20.470 ;
        RECT 75.860 19.675 76.120 19.935 ;
        RECT 76.180 19.675 76.440 19.935 ;
        RECT 76.500 19.675 76.760 19.935 ;
        RECT 94.095 20.235 94.355 20.495 ;
        RECT 94.765 20.235 95.025 20.495 ;
        RECT 97.045 20.235 97.305 20.495 ;
        RECT 99.325 20.235 99.585 20.495 ;
        RECT 101.605 20.235 101.865 20.495 ;
        RECT 103.885 20.235 104.145 20.495 ;
        RECT 106.165 20.235 106.425 20.495 ;
        RECT 108.445 20.235 108.705 20.495 ;
        RECT 110.725 20.235 110.985 20.495 ;
        RECT 113.005 20.235 113.265 20.495 ;
        RECT 115.285 20.235 115.545 20.495 ;
        RECT 117.565 20.235 117.825 20.495 ;
        RECT 118.235 20.235 118.495 20.495 ;
        RECT 99.760 19.630 100.020 19.890 ;
        RECT 100.080 19.630 100.340 19.890 ;
        RECT 100.400 19.630 100.660 19.890 ;
        RECT 101.605 18.695 101.865 18.955 ;
        RECT 101.605 18.375 101.865 18.635 ;
        RECT 55.935 16.525 56.195 16.785 ;
        RECT 56.605 16.525 56.865 16.785 ;
        RECT 57.385 16.525 57.645 16.785 ;
        RECT 58.165 16.525 58.425 16.785 ;
        RECT 60.445 16.525 60.705 16.785 ;
        RECT 62.725 16.525 62.985 16.785 ;
        RECT 63.505 16.525 63.765 16.785 ;
        RECT 64.285 16.525 64.545 16.785 ;
        RECT 64.955 16.525 65.215 16.785 ;
        RECT 60.125 15.920 60.385 16.180 ;
        RECT 60.445 15.920 60.705 16.180 ;
        RECT 60.765 15.920 61.025 16.180 ;
        RECT 72.810 17.130 73.070 17.390 ;
        RECT 73.130 17.130 73.390 17.390 ;
        RECT 73.450 17.130 73.710 17.390 ;
        RECT 69.145 16.525 69.405 16.785 ;
        RECT 69.815 16.525 70.075 16.785 ;
        RECT 71.095 16.525 71.355 16.785 ;
        RECT 72.375 16.525 72.635 16.785 ;
        RECT 76.935 16.525 77.195 16.785 ;
        RECT 78.215 16.525 78.475 16.785 ;
        RECT 79.495 16.525 79.755 16.785 ;
        RECT 80.775 16.525 81.035 16.785 ;
        RECT 82.055 16.525 82.315 16.785 ;
        RECT 84.335 16.525 84.595 16.785 ;
        RECT 86.615 16.525 86.875 16.785 ;
        RECT 87.895 16.525 88.155 16.785 ;
        RECT 89.175 16.525 89.435 16.785 ;
        RECT 89.845 16.525 90.105 16.785 ;
        RECT 72.675 15.920 72.935 16.180 ;
        RECT 72.995 15.920 73.255 16.180 ;
        RECT 73.315 15.920 73.575 16.180 ;
        RECT 84.015 15.915 84.275 16.175 ;
        RECT 84.335 15.915 84.595 16.175 ;
        RECT 84.655 15.915 84.915 16.175 ;
        RECT 101.605 18.055 101.865 18.315 ;
        RECT 106.165 18.695 106.425 18.955 ;
        RECT 106.165 18.375 106.425 18.635 ;
        RECT 137.035 21.350 137.295 21.610 ;
        RECT 135.075 20.870 135.335 21.130 ;
        RECT 135.075 20.550 135.335 20.810 ;
        RECT 135.075 20.230 135.335 20.490 ;
        RECT 135.745 20.870 136.005 21.130 ;
        RECT 135.745 20.550 136.005 20.810 ;
        RECT 135.745 20.230 136.005 20.490 ;
        RECT 136.175 20.870 136.435 21.130 ;
        RECT 136.175 20.550 136.435 20.810 ;
        RECT 136.175 20.230 136.435 20.490 ;
        RECT 136.605 20.870 136.865 21.130 ;
        RECT 136.605 20.550 136.865 20.810 ;
        RECT 136.605 20.230 136.865 20.490 ;
        RECT 137.035 21.030 137.295 21.290 ;
        RECT 137.895 21.350 138.155 21.610 ;
        RECT 137.035 20.710 137.295 20.970 ;
        RECT 137.035 20.390 137.295 20.650 ;
        RECT 137.035 20.070 137.295 20.330 ;
        RECT 137.465 20.870 137.725 21.130 ;
        RECT 137.465 20.550 137.725 20.810 ;
        RECT 137.465 20.230 137.725 20.490 ;
        RECT 137.895 21.030 138.155 21.290 ;
        RECT 138.755 21.350 139.015 21.610 ;
        RECT 137.895 20.710 138.155 20.970 ;
        RECT 137.895 20.390 138.155 20.650 ;
        RECT 137.035 19.750 137.295 20.010 ;
        RECT 137.895 20.070 138.155 20.330 ;
        RECT 138.325 20.870 138.585 21.130 ;
        RECT 138.325 20.550 138.585 20.810 ;
        RECT 138.325 20.230 138.585 20.490 ;
        RECT 138.755 21.030 139.015 21.290 ;
        RECT 139.615 21.350 139.875 21.610 ;
        RECT 138.755 20.710 139.015 20.970 ;
        RECT 138.755 20.390 139.015 20.650 ;
        RECT 137.895 19.750 138.155 20.010 ;
        RECT 138.755 20.070 139.015 20.330 ;
        RECT 139.185 20.870 139.445 21.130 ;
        RECT 139.185 20.550 139.445 20.810 ;
        RECT 139.185 20.230 139.445 20.490 ;
        RECT 139.615 21.030 139.875 21.290 ;
        RECT 140.475 21.350 140.735 21.610 ;
        RECT 139.615 20.710 139.875 20.970 ;
        RECT 139.615 20.390 139.875 20.650 ;
        RECT 138.755 19.750 139.015 20.010 ;
        RECT 139.615 20.070 139.875 20.330 ;
        RECT 140.045 20.870 140.305 21.130 ;
        RECT 140.045 20.550 140.305 20.810 ;
        RECT 140.045 20.230 140.305 20.490 ;
        RECT 140.475 21.030 140.735 21.290 ;
        RECT 141.335 21.350 141.595 21.610 ;
        RECT 140.475 20.710 140.735 20.970 ;
        RECT 140.475 20.390 140.735 20.650 ;
        RECT 139.615 19.750 139.875 20.010 ;
        RECT 140.475 20.070 140.735 20.330 ;
        RECT 140.905 20.870 141.165 21.130 ;
        RECT 140.905 20.550 141.165 20.810 ;
        RECT 140.905 20.230 141.165 20.490 ;
        RECT 141.335 21.030 141.595 21.290 ;
        RECT 142.195 21.350 142.455 21.610 ;
        RECT 141.335 20.710 141.595 20.970 ;
        RECT 141.335 20.390 141.595 20.650 ;
        RECT 140.475 19.750 140.735 20.010 ;
        RECT 141.335 20.070 141.595 20.330 ;
        RECT 141.765 20.870 142.025 21.130 ;
        RECT 141.765 20.550 142.025 20.810 ;
        RECT 141.765 20.230 142.025 20.490 ;
        RECT 142.195 21.030 142.455 21.290 ;
        RECT 142.195 20.710 142.455 20.970 ;
        RECT 142.195 20.390 142.455 20.650 ;
        RECT 141.335 19.750 141.595 20.010 ;
        RECT 142.195 20.070 142.455 20.330 ;
        RECT 142.625 20.870 142.885 21.130 ;
        RECT 142.625 20.550 142.885 20.810 ;
        RECT 142.625 20.230 142.885 20.490 ;
        RECT 143.055 20.870 143.315 21.130 ;
        RECT 143.055 20.550 143.315 20.810 ;
        RECT 143.055 20.230 143.315 20.490 ;
        RECT 143.485 20.870 143.745 21.130 ;
        RECT 143.485 20.550 143.745 20.810 ;
        RECT 143.485 20.230 143.745 20.490 ;
        RECT 144.155 20.870 144.415 21.130 ;
        RECT 144.155 20.550 144.415 20.810 ;
        RECT 144.155 20.230 144.415 20.490 ;
        RECT 142.195 19.750 142.455 20.010 ;
        RECT 135.840 18.375 136.100 18.635 ;
        RECT 136.160 18.375 136.420 18.635 ;
        RECT 106.165 18.055 106.425 18.315 ;
        RECT 99.760 16.540 100.020 16.800 ;
        RECT 100.080 16.540 100.340 16.800 ;
        RECT 100.400 16.540 100.660 16.800 ;
        RECT 94.095 16.005 94.355 16.265 ;
        RECT 94.095 15.685 94.355 15.945 ;
        RECT 94.095 15.365 94.355 15.625 ;
        RECT 94.765 16.005 95.025 16.265 ;
        RECT 94.765 15.685 95.025 15.945 ;
        RECT 94.765 15.365 95.025 15.625 ;
        RECT 97.045 16.005 97.305 16.265 ;
        RECT 97.045 15.685 97.305 15.945 ;
        RECT 97.045 15.365 97.305 15.625 ;
        RECT 99.325 16.005 99.585 16.265 ;
        RECT 99.325 15.685 99.585 15.945 ;
        RECT 99.325 15.365 99.585 15.625 ;
        RECT 101.605 16.005 101.865 16.265 ;
        RECT 101.605 15.685 101.865 15.945 ;
        RECT 101.605 15.365 101.865 15.625 ;
        RECT 103.885 16.005 104.145 16.265 ;
        RECT 103.885 15.685 104.145 15.945 ;
        RECT 103.885 15.365 104.145 15.625 ;
        RECT 106.165 16.005 106.425 16.265 ;
        RECT 106.165 15.685 106.425 15.945 ;
        RECT 106.165 15.365 106.425 15.625 ;
        RECT 108.445 16.005 108.705 16.265 ;
        RECT 108.445 15.685 108.705 15.945 ;
        RECT 108.445 15.365 108.705 15.625 ;
        RECT 110.725 16.005 110.985 16.265 ;
        RECT 110.725 15.685 110.985 15.945 ;
        RECT 110.725 15.365 110.985 15.625 ;
        RECT 113.005 16.005 113.265 16.265 ;
        RECT 113.005 15.685 113.265 15.945 ;
        RECT 113.005 15.365 113.265 15.625 ;
        RECT 115.285 16.005 115.545 16.265 ;
        RECT 115.285 15.685 115.545 15.945 ;
        RECT 115.285 15.365 115.545 15.625 ;
        RECT 117.565 16.005 117.825 16.265 ;
        RECT 117.565 15.685 117.825 15.945 ;
        RECT 117.565 15.365 117.825 15.625 ;
        RECT 118.235 16.005 118.495 16.265 ;
        RECT 118.235 15.685 118.495 15.945 ;
        RECT 137.895 18.695 138.155 18.955 ;
        RECT 137.895 18.375 138.155 18.635 ;
        RECT 137.895 18.055 138.155 18.315 ;
        RECT 135.075 17.020 135.335 17.280 ;
        RECT 135.075 16.700 135.335 16.960 ;
        RECT 135.075 16.380 135.335 16.640 ;
        RECT 135.745 17.020 136.005 17.280 ;
        RECT 135.745 16.700 136.005 16.960 ;
        RECT 135.745 16.380 136.005 16.640 ;
        RECT 136.175 17.020 136.435 17.280 ;
        RECT 136.175 16.700 136.435 16.960 ;
        RECT 136.175 16.380 136.435 16.640 ;
        RECT 136.605 17.020 136.865 17.280 ;
        RECT 136.605 16.700 136.865 16.960 ;
        RECT 136.605 16.380 136.865 16.640 ;
        RECT 137.035 17.020 137.295 17.280 ;
        RECT 137.035 16.700 137.295 16.960 ;
        RECT 137.035 16.380 137.295 16.640 ;
        RECT 137.465 17.020 137.725 17.280 ;
        RECT 137.465 16.700 137.725 16.960 ;
        RECT 137.465 16.380 137.725 16.640 ;
        RECT 137.895 17.020 138.155 17.280 ;
        RECT 137.895 16.700 138.155 16.960 ;
        RECT 137.895 16.380 138.155 16.640 ;
        RECT 138.325 17.020 138.585 17.280 ;
        RECT 138.325 16.700 138.585 16.960 ;
        RECT 138.325 16.380 138.585 16.640 ;
        RECT 138.755 17.020 139.015 17.280 ;
        RECT 138.755 16.700 139.015 16.960 ;
        RECT 138.755 16.380 139.015 16.640 ;
        RECT 139.185 17.020 139.445 17.280 ;
        RECT 139.185 16.700 139.445 16.960 ;
        RECT 139.185 16.380 139.445 16.640 ;
        RECT 139.615 17.020 139.875 17.280 ;
        RECT 139.615 16.700 139.875 16.960 ;
        RECT 139.615 16.380 139.875 16.640 ;
        RECT 140.045 17.020 140.305 17.280 ;
        RECT 140.045 16.700 140.305 16.960 ;
        RECT 140.045 16.380 140.305 16.640 ;
        RECT 140.475 17.020 140.735 17.280 ;
        RECT 140.475 16.700 140.735 16.960 ;
        RECT 140.475 16.380 140.735 16.640 ;
        RECT 140.905 17.020 141.165 17.280 ;
        RECT 140.905 16.700 141.165 16.960 ;
        RECT 140.905 16.380 141.165 16.640 ;
        RECT 141.335 17.020 141.595 17.280 ;
        RECT 141.335 16.700 141.595 16.960 ;
        RECT 141.335 16.380 141.595 16.640 ;
        RECT 141.765 17.020 142.025 17.280 ;
        RECT 141.765 16.700 142.025 16.960 ;
        RECT 141.765 16.380 142.025 16.640 ;
        RECT 142.195 17.020 142.455 17.280 ;
        RECT 142.195 16.700 142.455 16.960 ;
        RECT 142.195 16.380 142.455 16.640 ;
        RECT 142.625 17.020 142.885 17.280 ;
        RECT 142.625 16.700 142.885 16.960 ;
        RECT 142.625 16.380 142.885 16.640 ;
        RECT 143.055 17.020 143.315 17.280 ;
        RECT 143.055 16.700 143.315 16.960 ;
        RECT 143.055 16.380 143.315 16.640 ;
        RECT 143.485 17.020 143.745 17.280 ;
        RECT 143.485 16.700 143.745 16.960 ;
        RECT 143.485 16.380 143.745 16.640 ;
        RECT 144.155 17.020 144.415 17.280 ;
        RECT 144.155 16.700 144.415 16.960 ;
        RECT 144.155 16.380 144.415 16.640 ;
        RECT 118.235 15.365 118.495 15.625 ;
        RECT 58.600 12.965 58.860 13.225 ;
        RECT 58.920 12.965 59.180 13.225 ;
        RECT 59.240 12.965 59.500 13.225 ;
        RECT 66.280 12.965 66.540 13.225 ;
        RECT 66.600 12.965 66.860 13.225 ;
        RECT 66.920 12.965 67.180 13.225 ;
        RECT 92.130 12.965 92.390 13.225 ;
        RECT 92.450 12.965 92.710 13.225 ;
        RECT 92.770 12.965 93.030 13.225 ;
        RECT 55.935 12.430 56.195 12.690 ;
        RECT 55.935 12.110 56.195 12.370 ;
        RECT 55.935 11.790 56.195 12.050 ;
        RECT 56.605 12.430 56.865 12.690 ;
        RECT 56.605 12.110 56.865 12.370 ;
        RECT 56.605 11.790 56.865 12.050 ;
        RECT 57.385 12.430 57.645 12.690 ;
        RECT 57.385 12.110 57.645 12.370 ;
        RECT 57.385 11.790 57.645 12.050 ;
        RECT 58.165 12.430 58.425 12.690 ;
        RECT 58.165 12.110 58.425 12.370 ;
        RECT 58.165 11.790 58.425 12.050 ;
        RECT 60.445 12.430 60.705 12.690 ;
        RECT 60.445 12.110 60.705 12.370 ;
        RECT 60.445 11.790 60.705 12.050 ;
        RECT 62.725 12.430 62.985 12.690 ;
        RECT 62.725 12.110 62.985 12.370 ;
        RECT 62.725 11.790 62.985 12.050 ;
        RECT 63.505 12.430 63.765 12.690 ;
        RECT 63.505 12.110 63.765 12.370 ;
        RECT 63.505 11.790 63.765 12.050 ;
        RECT 64.285 12.430 64.545 12.690 ;
        RECT 64.285 12.110 64.545 12.370 ;
        RECT 64.285 11.790 64.545 12.050 ;
        RECT 65.065 12.430 65.325 12.690 ;
        RECT 65.065 12.110 65.325 12.370 ;
        RECT 65.065 11.790 65.325 12.050 ;
        RECT 65.845 12.430 66.105 12.690 ;
        RECT 65.845 12.110 66.105 12.370 ;
        RECT 65.845 11.790 66.105 12.050 ;
        RECT 68.125 12.430 68.385 12.690 ;
        RECT 68.125 12.110 68.385 12.370 ;
        RECT 68.125 11.790 68.385 12.050 ;
        RECT 70.405 12.430 70.665 12.690 ;
        RECT 70.405 12.110 70.665 12.370 ;
        RECT 70.405 11.790 70.665 12.050 ;
        RECT 72.685 12.430 72.945 12.690 ;
        RECT 72.685 12.110 72.945 12.370 ;
        RECT 72.685 11.790 72.945 12.050 ;
        RECT 74.965 12.430 75.225 12.690 ;
        RECT 74.965 12.110 75.225 12.370 ;
        RECT 74.965 11.790 75.225 12.050 ;
        RECT 77.245 12.430 77.505 12.690 ;
        RECT 77.245 12.110 77.505 12.370 ;
        RECT 77.245 11.790 77.505 12.050 ;
        RECT 79.525 12.430 79.785 12.690 ;
        RECT 79.525 12.110 79.785 12.370 ;
        RECT 79.525 11.790 79.785 12.050 ;
        RECT 81.805 12.430 82.065 12.690 ;
        RECT 81.805 12.110 82.065 12.370 ;
        RECT 81.805 11.790 82.065 12.050 ;
        RECT 84.085 12.430 84.345 12.690 ;
        RECT 84.085 12.110 84.345 12.370 ;
        RECT 84.085 11.790 84.345 12.050 ;
        RECT 86.365 12.430 86.625 12.690 ;
        RECT 86.365 12.110 86.625 12.370 ;
        RECT 86.365 11.790 86.625 12.050 ;
        RECT 88.645 12.430 88.905 12.690 ;
        RECT 88.645 12.110 88.905 12.370 ;
        RECT 88.645 11.790 88.905 12.050 ;
        RECT 90.925 12.430 91.185 12.690 ;
        RECT 90.925 12.110 91.185 12.370 ;
        RECT 90.925 11.790 91.185 12.050 ;
        RECT 93.205 12.430 93.465 12.690 ;
        RECT 93.205 12.110 93.465 12.370 ;
        RECT 93.205 11.790 93.465 12.050 ;
        RECT 93.985 12.430 94.245 12.690 ;
        RECT 93.985 12.110 94.245 12.370 ;
        RECT 93.985 11.790 94.245 12.050 ;
        RECT 94.765 12.430 95.025 12.690 ;
        RECT 94.765 12.110 95.025 12.370 ;
        RECT 94.765 11.790 95.025 12.050 ;
        RECT 95.435 12.430 95.695 12.690 ;
        RECT 95.435 12.110 95.695 12.370 ;
        RECT 95.435 11.790 95.695 12.050 ;
        RECT 55.935 8.840 56.195 9.100 ;
        RECT 55.935 8.520 56.195 8.780 ;
        RECT 55.935 8.200 56.195 8.460 ;
        RECT 65.845 8.840 66.105 9.100 ;
        RECT 65.845 8.520 66.105 8.780 ;
        RECT 65.845 8.200 66.105 8.460 ;
        RECT 68.125 8.840 68.385 9.100 ;
        RECT 68.125 8.520 68.385 8.780 ;
        RECT 68.125 8.200 68.385 8.460 ;
        RECT 70.405 8.840 70.665 9.100 ;
        RECT 70.405 8.520 70.665 8.780 ;
        RECT 70.405 8.200 70.665 8.460 ;
        RECT 72.685 8.840 72.945 9.100 ;
        RECT 72.685 8.520 72.945 8.780 ;
        RECT 72.685 8.200 72.945 8.460 ;
        RECT 74.965 8.840 75.225 9.100 ;
        RECT 74.965 8.520 75.225 8.780 ;
        RECT 74.965 8.200 75.225 8.460 ;
        RECT 77.245 8.840 77.505 9.100 ;
        RECT 77.245 8.520 77.505 8.780 ;
        RECT 77.245 8.200 77.505 8.460 ;
        RECT 79.525 8.840 79.785 9.100 ;
        RECT 79.525 8.520 79.785 8.780 ;
        RECT 79.525 8.200 79.785 8.460 ;
        RECT 81.805 8.840 82.065 9.100 ;
        RECT 81.805 8.520 82.065 8.780 ;
        RECT 81.805 8.200 82.065 8.460 ;
        RECT 84.085 8.840 84.345 9.100 ;
        RECT 84.085 8.520 84.345 8.780 ;
        RECT 84.085 8.200 84.345 8.460 ;
        RECT 86.365 8.840 86.625 9.100 ;
        RECT 86.365 8.520 86.625 8.780 ;
        RECT 86.365 8.200 86.625 8.460 ;
        RECT 88.645 8.840 88.905 9.100 ;
        RECT 88.645 8.520 88.905 8.780 ;
        RECT 88.645 8.200 88.905 8.460 ;
        RECT 90.925 8.840 91.185 9.100 ;
        RECT 90.925 8.520 91.185 8.780 ;
        RECT 90.925 8.200 91.185 8.460 ;
        RECT 93.205 8.840 93.465 9.100 ;
        RECT 93.205 8.520 93.465 8.780 ;
        RECT 93.205 8.200 93.465 8.460 ;
        RECT 95.435 8.840 95.695 9.100 ;
        RECT 95.435 8.520 95.695 8.780 ;
        RECT 95.435 8.200 95.695 8.460 ;
        RECT 79.205 7.665 79.465 7.925 ;
        RECT 79.525 7.665 79.785 7.925 ;
        RECT 79.845 7.665 80.105 7.925 ;
      LAYER met2 ;
        RECT -4.050 108.665 -2.970 109.265 ;
        RECT 202.090 108.665 203.570 109.265 ;
        RECT -4.880 78.375 -4.550 95.155 ;
        RECT -4.050 66.355 -3.720 108.665 ;
        RECT -2.390 107.565 -1.710 108.165 ;
        RECT -3.220 71.335 -2.890 98.830 ;
        RECT -2.390 74.680 -1.790 107.565 ;
        RECT -1.290 68.715 -0.690 93.530 ;
        RECT 141.615 78.395 142.785 78.725 ;
        RECT 142.035 77.625 142.365 78.395 ;
        RECT 141.750 77.305 142.650 77.625 ;
        RECT 137.110 76.425 137.400 77.125 ;
        RECT 137.745 76.425 138.025 77.125 ;
        RECT 138.175 76.425 138.455 77.125 ;
        RECT 138.605 76.425 138.885 77.125 ;
        RECT 139.035 76.425 139.315 77.125 ;
        RECT 139.465 76.425 139.745 77.125 ;
        RECT 139.895 76.425 140.175 77.125 ;
        RECT 140.325 76.425 140.605 77.125 ;
        RECT 140.755 76.425 141.035 77.125 ;
        RECT 141.185 76.425 141.465 77.125 ;
        RECT 141.615 76.240 141.895 77.125 ;
        RECT 142.045 76.425 142.325 77.125 ;
        RECT 142.475 76.240 142.755 77.125 ;
        RECT 142.905 76.425 143.185 77.125 ;
        RECT 143.335 76.425 143.615 77.125 ;
        RECT 143.765 76.425 144.045 77.125 ;
        RECT 144.195 76.425 144.475 77.125 ;
        RECT 144.625 76.425 144.905 77.125 ;
        RECT 145.055 76.425 145.335 77.125 ;
        RECT 145.485 76.425 145.765 77.125 ;
        RECT 145.915 76.425 146.195 77.125 ;
        RECT 146.345 76.425 146.625 77.125 ;
        RECT 146.970 76.425 147.260 77.125 ;
        RECT 42.710 75.180 43.000 75.880 ;
        RECT 43.345 75.180 43.625 75.880 ;
        RECT 45.625 75.180 45.905 75.880 ;
        RECT 47.905 75.010 48.185 75.880 ;
        RECT 50.185 75.180 50.465 75.880 ;
        RECT 52.465 75.010 52.745 75.880 ;
        RECT 54.745 75.180 55.025 75.880 ;
        RECT 57.025 75.010 57.305 75.880 ;
        RECT 59.305 75.180 59.585 75.880 ;
        RECT 61.585 75.010 61.865 75.880 ;
        RECT 63.865 75.180 64.145 75.880 ;
        RECT 66.145 75.010 66.425 75.880 ;
        RECT 68.425 75.180 68.705 75.880 ;
        RECT 70.705 75.010 70.985 75.880 ;
        RECT 72.985 75.180 73.265 75.880 ;
        RECT 75.265 75.010 75.545 75.880 ;
        RECT 77.545 75.180 77.825 75.880 ;
        RECT 79.825 75.010 80.105 75.880 ;
        RECT 82.105 75.180 82.385 75.880 ;
        RECT 41.070 74.680 80.105 75.010 ;
        RECT 42.710 73.810 43.000 74.510 ;
        RECT 43.345 73.810 43.625 74.510 ;
        RECT 45.625 73.810 45.905 74.510 ;
        RECT 47.905 73.810 48.185 74.680 ;
        RECT 50.185 73.810 50.465 74.510 ;
        RECT 52.465 73.810 52.745 74.680 ;
        RECT 54.745 73.810 55.025 74.510 ;
        RECT 57.025 73.810 57.305 74.680 ;
        RECT 59.305 73.810 59.585 74.510 ;
        RECT 61.585 73.810 61.865 74.680 ;
        RECT 63.865 73.810 64.145 74.510 ;
        RECT 66.145 73.810 66.425 74.680 ;
        RECT 68.425 73.810 68.705 74.510 ;
        RECT 70.705 73.810 70.985 74.680 ;
        RECT 72.985 73.810 73.265 74.510 ;
        RECT 75.265 73.810 75.545 74.680 ;
        RECT 77.545 73.810 77.825 74.510 ;
        RECT 79.825 73.810 80.105 74.680 ;
        RECT 82.105 73.810 82.385 74.510 ;
        RECT 84.385 73.065 84.665 75.880 ;
        RECT 86.665 75.180 86.945 75.880 ;
        RECT 86.665 73.810 86.945 74.510 ;
        RECT 88.945 73.065 89.225 75.880 ;
        RECT 91.225 75.180 91.505 75.880 ;
        RECT 91.225 73.810 91.505 74.510 ;
        RECT 93.505 73.065 93.785 75.880 ;
        RECT 95.785 75.180 96.065 75.880 ;
        RECT 95.785 73.810 96.065 74.510 ;
        RECT 98.065 73.065 98.345 75.880 ;
        RECT 100.345 75.180 100.625 75.880 ;
        RECT 100.345 73.810 100.625 74.510 ;
        RECT 102.625 73.065 102.905 75.880 ;
        RECT 104.905 75.180 105.185 75.880 ;
        RECT 104.905 73.810 105.185 74.510 ;
        RECT 107.185 73.065 107.465 75.880 ;
        RECT 109.465 75.180 109.745 75.880 ;
        RECT 109.465 73.810 109.745 74.510 ;
        RECT 111.745 73.065 112.025 75.880 ;
        RECT 114.025 75.180 114.305 75.880 ;
        RECT 114.025 73.810 114.305 74.510 ;
        RECT 116.305 73.065 116.585 75.880 ;
        RECT 118.585 75.180 118.865 75.880 ;
        RECT 120.865 75.180 121.145 75.880 ;
        RECT 123.145 75.180 123.425 75.880 ;
        RECT 125.425 75.180 125.705 75.880 ;
        RECT 127.705 75.180 127.985 75.880 ;
        RECT 129.985 75.180 130.265 75.880 ;
        RECT 130.610 75.180 130.900 75.880 ;
        RECT 141.615 75.640 152.135 76.240 ;
        RECT 168.605 75.640 169.205 93.530 ;
        RECT 185.955 75.640 187.035 76.240 ;
        RECT 141.615 75.290 141.895 75.640 ;
        RECT 142.475 75.290 142.755 75.640 ;
        RECT 123.980 74.680 124.880 75.010 ;
        RECT 136.120 74.960 137.290 75.290 ;
        RECT 139.035 74.960 145.425 75.290 ;
        RECT 118.585 73.810 118.865 74.510 ;
        RECT 120.865 73.810 121.145 74.510 ;
        RECT 123.145 73.810 123.425 74.510 ;
        RECT 124.290 73.620 124.570 74.680 ;
        RECT 123.950 73.330 124.910 73.620 ;
        RECT 84.385 72.785 116.585 73.065 ;
        RECT 93.125 71.355 94.295 71.685 ;
        RECT 0.605 68.695 1.685 69.065 ;
        RECT 93.145 69.045 93.425 71.165 ;
        RECT 94.005 69.045 94.285 71.165 ;
        RECT 90.760 68.715 96.570 69.045 ;
        RECT 0.605 57.100 1.205 68.695 ;
        RECT 39.625 67.785 40.795 68.115 ;
        RECT 33.520 63.045 33.810 64.045 ;
        RECT 34.195 63.045 34.475 64.045 ;
        RECT 34.625 63.045 34.905 64.045 ;
        RECT 35.055 63.045 35.335 64.045 ;
        RECT 35.485 61.535 35.765 64.545 ;
        RECT 35.915 63.045 36.195 64.045 ;
        RECT 36.345 61.535 36.625 64.545 ;
        RECT 36.775 63.045 37.055 64.045 ;
        RECT 37.205 63.045 37.485 64.045 ;
        RECT 37.635 63.045 37.915 64.045 ;
        RECT 38.300 63.045 38.590 64.045 ;
        RECT 34.205 61.205 34.975 61.535 ;
        RECT 35.485 61.525 37.860 61.535 ;
        RECT 40.045 61.525 40.375 67.785 ;
        RECT 90.760 66.895 91.040 68.715 ;
        RECT 90.220 66.375 90.990 66.705 ;
        RECT 91.190 65.615 91.470 67.595 ;
        RECT 91.620 66.895 91.900 68.715 ;
        RECT 95.430 66.895 95.710 68.715 ;
        RECT 95.860 65.615 96.140 67.595 ;
        RECT 96.290 66.895 96.570 68.715 ;
        RECT 96.770 67.785 97.540 68.115 ;
        RECT 72.985 65.285 107.560 65.615 ;
        RECT 42.670 63.345 42.960 64.045 ;
        RECT 43.345 63.345 43.625 64.045 ;
        RECT 45.625 63.345 45.905 64.045 ;
        RECT 47.905 63.345 48.185 64.045 ;
        RECT 50.185 63.175 50.465 64.045 ;
        RECT 52.465 63.345 52.745 64.045 ;
        RECT 54.745 63.175 55.025 64.045 ;
        RECT 57.025 63.345 57.305 64.045 ;
        RECT 59.305 63.175 59.585 64.045 ;
        RECT 61.585 63.345 61.865 64.045 ;
        RECT 63.865 63.175 64.145 64.045 ;
        RECT 66.145 63.345 66.425 64.045 ;
        RECT 68.425 63.175 68.705 64.045 ;
        RECT 70.705 63.345 70.985 64.045 ;
        RECT 50.185 62.845 68.705 63.175 ;
        RECT 42.670 61.975 42.960 62.675 ;
        RECT 43.345 61.975 43.625 62.675 ;
        RECT 45.625 61.975 45.905 62.675 ;
        RECT 47.905 61.975 48.185 62.675 ;
        RECT 35.485 61.205 40.375 61.525 ;
        RECT 50.185 61.805 50.465 62.845 ;
        RECT 52.465 61.975 52.745 62.675 ;
        RECT 54.745 61.805 55.025 62.845 ;
        RECT 57.025 61.975 57.305 62.675 ;
        RECT 59.305 61.805 59.585 62.845 ;
        RECT 61.585 61.975 61.865 62.675 ;
        RECT 63.865 61.805 64.145 62.845 ;
        RECT 66.145 61.975 66.425 62.675 ;
        RECT 68.425 61.805 68.705 62.845 ;
        RECT 70.705 61.975 70.985 62.675 ;
        RECT 50.185 61.475 68.705 61.805 ;
        RECT 33.520 59.195 33.810 60.195 ;
        RECT 34.195 59.195 34.475 60.195 ;
        RECT 34.625 59.195 34.905 60.195 ;
        RECT 35.055 59.195 35.335 60.195 ;
        RECT 35.485 59.195 35.765 61.205 ;
        RECT 35.915 59.195 36.195 60.195 ;
        RECT 36.345 59.195 36.625 61.205 ;
        RECT 36.980 61.195 40.375 61.205 ;
        RECT 42.670 60.605 42.960 61.305 ;
        RECT 43.345 60.605 43.625 61.305 ;
        RECT 45.625 60.605 45.905 61.305 ;
        RECT 47.905 60.605 48.185 61.305 ;
        RECT 50.185 60.605 50.465 61.475 ;
        RECT 52.465 60.605 52.745 61.305 ;
        RECT 54.745 60.605 55.025 61.475 ;
        RECT 57.025 60.605 57.305 61.305 ;
        RECT 59.305 60.605 59.585 61.475 ;
        RECT 61.585 60.605 61.865 61.305 ;
        RECT 63.865 60.605 64.145 61.475 ;
        RECT 66.145 60.605 66.425 61.305 ;
        RECT 68.425 60.605 68.705 61.475 ;
        RECT 70.705 60.605 70.985 61.305 ;
        RECT 72.985 60.605 73.265 65.285 ;
        RECT 75.265 63.345 75.545 64.045 ;
        RECT 75.265 61.975 75.545 62.675 ;
        RECT 75.265 60.605 75.545 61.305 ;
        RECT 77.545 60.605 77.825 65.285 ;
        RECT 79.825 63.345 80.105 64.045 ;
        RECT 79.825 61.975 80.105 62.675 ;
        RECT 79.825 60.605 80.105 61.305 ;
        RECT 82.105 60.605 82.385 65.285 ;
        RECT 84.385 63.345 84.665 64.045 ;
        RECT 84.385 61.975 84.665 62.675 ;
        RECT 84.385 60.605 84.665 61.305 ;
        RECT 86.665 60.605 86.945 65.285 ;
        RECT 88.945 63.345 89.225 64.045 ;
        RECT 88.945 61.975 89.225 62.675 ;
        RECT 88.945 60.605 89.225 61.305 ;
        RECT 91.225 60.605 91.505 65.285 ;
        RECT 93.505 63.345 93.785 64.045 ;
        RECT 93.505 61.975 93.785 62.675 ;
        RECT 93.505 60.605 93.785 61.305 ;
        RECT 95.785 60.605 96.065 65.285 ;
        RECT 98.065 63.345 98.345 64.045 ;
        RECT 98.065 61.975 98.345 62.675 ;
        RECT 98.065 60.605 98.345 61.305 ;
        RECT 100.345 60.605 100.625 65.285 ;
        RECT 102.625 63.345 102.905 64.045 ;
        RECT 102.625 61.975 102.905 62.675 ;
        RECT 102.625 60.605 102.905 61.305 ;
        RECT 104.905 60.605 105.185 65.285 ;
        RECT 107.185 63.345 107.465 64.045 ;
        RECT 108.255 63.175 108.755 72.785 ;
        RECT 125.425 72.485 125.705 74.510 ;
        RECT 127.705 73.810 127.985 74.510 ;
        RECT 129.985 73.810 130.265 74.510 ;
        RECT 130.610 73.810 130.900 74.510 ;
        RECT 125.425 72.155 126.595 72.485 ;
        RECT 127.325 71.355 128.495 71.685 ;
        RECT 136.120 71.660 136.450 74.960 ;
        RECT 137.595 74.045 138.630 74.375 ;
        RECT 138.605 72.155 138.885 73.855 ;
        RECT 136.120 71.330 138.250 71.660 ;
        RECT 127.345 69.045 127.625 71.165 ;
        RECT 128.205 69.045 128.485 71.165 ;
        RECT 139.035 71.140 139.315 74.960 ;
        RECT 139.465 72.155 139.745 73.855 ;
        RECT 139.895 71.140 140.175 74.960 ;
        RECT 140.325 72.155 140.605 73.855 ;
        RECT 143.855 72.155 144.135 73.855 ;
        RECT 142.935 71.440 144.025 71.770 ;
        RECT 144.285 71.140 144.565 74.960 ;
        RECT 144.715 72.155 144.995 73.855 ;
        RECT 145.145 71.140 145.425 74.960 ;
        RECT 145.920 74.940 146.600 75.310 ;
        RECT 146.095 74.375 146.425 74.940 ;
        RECT 145.970 74.045 146.550 74.375 ;
        RECT 145.575 72.135 145.855 73.855 ;
        RECT 147.920 71.420 148.250 74.395 ;
        RECT 137.070 70.440 137.360 71.140 ;
        RECT 137.745 70.440 138.025 71.140 ;
        RECT 138.175 70.440 138.455 71.140 ;
        RECT 138.605 69.045 138.885 71.140 ;
        RECT 139.030 70.440 139.315 71.140 ;
        RECT 139.465 69.045 139.745 71.140 ;
        RECT 139.890 70.440 140.175 71.140 ;
        RECT 140.325 69.045 140.605 71.140 ;
        RECT 140.755 70.440 141.035 71.140 ;
        RECT 141.185 70.440 141.465 71.140 ;
        RECT 142.995 70.440 143.275 71.140 ;
        RECT 143.425 70.440 143.705 71.140 ;
        RECT 143.855 69.045 144.135 71.140 ;
        RECT 144.280 70.440 144.565 71.140 ;
        RECT 144.715 69.045 144.995 71.140 ;
        RECT 145.140 70.440 145.425 71.140 ;
        RECT 145.575 69.045 145.855 71.140 ;
        RECT 146.005 70.440 146.285 71.140 ;
        RECT 146.435 70.440 146.715 71.140 ;
        RECT 147.060 70.440 147.350 71.140 ;
        RECT 124.960 68.715 130.770 69.045 ;
        RECT 138.605 68.715 145.855 69.045 ;
        RECT 124.960 66.895 125.240 68.715 ;
        RECT 124.420 66.375 125.190 66.705 ;
        RECT 125.390 65.615 125.670 67.595 ;
        RECT 125.820 66.895 126.100 68.715 ;
        RECT 129.630 66.895 129.910 68.715 ;
        RECT 130.060 65.615 130.340 67.595 ;
        RECT 130.490 66.895 130.770 68.715 ;
        RECT 130.970 67.785 131.740 68.115 ;
        RECT 132.015 66.745 132.305 67.445 ;
        RECT 136.790 66.745 137.080 67.445 ;
        RECT 137.465 66.745 137.745 67.445 ;
        RECT 139.745 66.745 140.025 67.445 ;
        RECT 142.025 66.745 142.305 68.715 ;
        RECT 144.305 66.745 144.585 67.445 ;
        RECT 146.585 66.745 146.865 67.445 ;
        RECT 147.250 66.745 147.540 67.445 ;
        RECT 137.960 66.225 138.860 66.555 ;
        RECT 109.465 65.285 114.305 65.615 ;
        RECT 107.895 62.845 109.115 63.175 ;
        RECT 107.185 61.975 107.465 62.675 ;
        RECT 107.185 60.605 107.465 61.305 ;
        RECT 109.465 60.605 109.745 65.285 ;
        RECT 111.745 63.345 112.025 64.045 ;
        RECT 111.745 61.975 112.025 62.675 ;
        RECT 111.745 60.605 112.025 61.305 ;
        RECT 114.025 60.605 114.305 65.285 ;
        RECT 118.585 65.285 137.105 65.615 ;
        RECT 116.305 63.345 116.585 64.045 ;
        RECT 116.305 61.975 116.585 62.675 ;
        RECT 116.305 60.605 116.585 61.305 ;
        RECT 118.585 60.605 118.865 65.285 ;
        RECT 120.865 63.345 121.145 64.045 ;
        RECT 120.865 61.975 121.145 62.675 ;
        RECT 120.865 60.605 121.145 61.305 ;
        RECT 123.145 60.605 123.425 65.285 ;
        RECT 125.425 63.345 125.705 64.045 ;
        RECT 125.425 61.975 125.705 62.675 ;
        RECT 125.425 60.605 125.705 61.305 ;
        RECT 127.705 60.605 127.985 65.285 ;
        RECT 129.985 63.345 130.265 64.045 ;
        RECT 129.985 61.975 130.265 62.675 ;
        RECT 129.985 60.605 130.265 61.305 ;
        RECT 132.265 60.605 132.545 65.285 ;
        RECT 134.545 63.345 134.825 64.045 ;
        RECT 134.545 61.975 134.825 62.675 ;
        RECT 134.545 60.605 134.825 61.305 ;
        RECT 136.825 60.605 137.105 65.285 ;
        RECT 137.960 63.175 138.240 66.225 ;
        RECT 139.105 63.345 139.385 64.045 ;
        RECT 141.385 63.345 141.665 64.045 ;
        RECT 143.665 63.345 143.945 64.045 ;
        RECT 144.330 63.345 144.620 64.045 ;
        RECT 137.650 62.845 138.550 63.175 ;
        RECT 139.105 61.975 139.385 62.675 ;
        RECT 141.385 61.975 141.665 62.675 ;
        RECT 143.665 61.975 143.945 62.675 ;
        RECT 144.330 61.975 144.620 62.675 ;
        RECT 139.105 60.605 139.385 61.305 ;
        RECT 141.385 60.605 141.665 61.305 ;
        RECT 143.665 60.605 143.945 61.305 ;
        RECT 144.330 60.605 144.620 61.305 ;
        RECT 36.775 59.195 37.055 60.195 ;
        RECT 37.205 59.195 37.485 60.195 ;
        RECT 37.635 59.195 37.915 60.195 ;
        RECT 38.300 59.195 38.590 60.195 ;
        RECT 33.855 39.630 35.025 39.930 ;
        RECT 32.755 35.950 33.925 36.250 ;
        RECT 33.325 -2.405 33.925 35.950 ;
        RECT 34.425 -1.305 35.025 39.630 ;
        RECT 52.850 29.045 53.450 57.700 ;
        RECT 53.950 57.100 55.030 57.700 ;
        RECT 53.950 29.045 54.550 57.100 ;
        RECT 186.195 55.670 186.795 75.640 ;
        RECT 120.560 55.070 121.640 55.670 ;
        RECT 185.690 55.070 186.795 55.670 ;
        RECT 187.345 74.960 188.515 75.290 ;
        RECT 78.650 53.360 79.820 53.690 ;
        RECT 79.490 53.160 79.820 53.360 ;
        RECT 79.205 52.830 80.105 53.160 ;
        RECT 55.920 51.640 56.210 52.640 ;
        RECT 65.835 51.640 66.115 52.640 ;
        RECT 68.115 51.640 68.395 52.640 ;
        RECT 70.395 51.640 70.675 52.640 ;
        RECT 72.675 51.640 72.955 52.640 ;
        RECT 74.955 51.640 75.235 52.640 ;
        RECT 77.235 51.640 77.515 52.640 ;
        RECT 79.515 50.535 79.795 52.640 ;
        RECT 81.795 51.640 82.075 52.640 ;
        RECT 84.075 51.640 84.355 52.640 ;
        RECT 86.355 51.640 86.635 52.640 ;
        RECT 88.635 51.640 88.915 52.640 ;
        RECT 90.915 51.640 91.195 52.640 ;
        RECT 93.195 51.640 93.475 52.640 ;
        RECT 95.420 51.640 95.710 52.640 ;
        RECT 65.835 50.205 93.475 50.535 ;
        RECT 55.920 48.050 56.210 49.050 ;
        RECT 56.595 48.050 56.875 49.050 ;
        RECT 57.375 48.050 57.655 49.050 ;
        RECT 58.155 48.050 58.435 49.050 ;
        RECT 58.600 47.530 59.500 47.860 ;
        RECT 55.440 38.480 55.720 46.640 ;
        RECT 58.600 46.620 58.890 47.530 ;
        RECT 57.720 46.290 58.890 46.620 ;
        RECT 60.435 46.355 60.715 49.050 ;
        RECT 62.715 48.050 62.995 49.050 ;
        RECT 63.495 48.050 63.775 49.050 ;
        RECT 64.275 48.050 64.555 49.050 ;
        RECT 65.055 48.050 65.335 49.050 ;
        RECT 65.835 48.050 66.115 50.205 ;
        RECT 66.280 47.530 67.180 47.860 ;
        RECT 60.435 45.695 61.605 46.025 ;
        RECT 60.435 44.905 60.715 45.695 ;
        RECT 60.125 44.575 61.025 44.905 ;
        RECT 55.920 43.885 56.210 44.385 ;
        RECT 56.595 43.885 56.875 44.385 ;
        RECT 57.375 43.885 57.655 44.385 ;
        RECT 58.155 43.885 58.435 44.385 ;
        RECT 55.440 38.150 56.610 38.480 ;
        RECT 60.435 37.655 60.715 44.385 ;
        RECT 62.715 43.885 62.995 44.385 ;
        RECT 63.495 43.885 63.775 44.385 ;
        RECT 64.275 43.885 64.555 44.385 ;
        RECT 64.940 43.885 65.230 44.385 ;
        RECT 60.435 37.325 61.605 37.655 ;
        RECT 66.280 36.750 66.610 47.530 ;
        RECT 68.115 46.355 68.395 49.050 ;
        RECT 70.395 48.050 70.675 50.205 ;
        RECT 72.675 44.905 72.955 49.050 ;
        RECT 74.955 48.050 75.235 50.205 ;
        RECT 77.235 46.355 77.515 49.050 ;
        RECT 79.515 48.050 79.795 50.205 ;
        RECT 81.795 46.355 82.075 49.050 ;
        RECT 84.075 48.050 84.355 50.205 ;
        RECT 83.880 46.375 85.050 46.705 ;
        RECT 84.325 46.025 84.605 46.375 ;
        RECT 86.355 46.355 86.635 49.050 ;
        RECT 88.635 48.050 88.915 50.205 ;
        RECT 90.915 46.355 91.195 49.050 ;
        RECT 93.195 48.050 93.475 50.205 ;
        RECT 93.975 48.050 94.255 49.050 ;
        RECT 94.755 48.050 95.035 49.050 ;
        RECT 95.420 48.050 95.710 49.050 ;
        RECT 92.130 47.530 93.030 47.860 ;
        RECT 83.435 45.695 84.605 46.025 ;
        RECT 84.325 44.910 84.605 45.695 ;
        RECT 72.675 44.575 73.575 44.905 ;
        RECT 84.015 44.580 84.915 44.910 ;
        RECT 69.130 43.885 69.420 44.385 ;
        RECT 69.805 43.885 70.085 44.385 ;
        RECT 71.085 43.885 71.365 44.385 ;
        RECT 72.365 43.885 72.645 44.385 ;
        RECT 76.925 43.885 77.205 44.385 ;
        RECT 78.205 43.885 78.485 44.385 ;
        RECT 79.485 43.885 79.765 44.385 ;
        RECT 80.765 43.885 81.045 44.385 ;
        RECT 82.045 43.885 82.325 44.385 ;
        RECT 84.325 43.885 84.605 44.580 ;
        RECT 86.605 43.885 86.885 44.385 ;
        RECT 87.885 43.885 88.165 44.385 ;
        RECT 89.165 43.885 89.445 44.385 ;
        RECT 89.830 43.885 90.120 44.385 ;
        RECT 72.810 43.365 73.710 43.695 ;
        RECT 73.120 42.110 73.400 43.365 ;
        RECT 75.280 42.460 76.450 42.790 ;
        RECT 73.120 41.780 74.290 42.110 ;
        RECT 76.170 41.150 76.450 42.460 ;
        RECT 75.860 40.820 76.760 41.150 ;
        RECT 69.130 39.630 69.420 40.630 ;
        RECT 69.805 39.630 70.085 40.630 ;
        RECT 71.085 39.630 71.365 40.630 ;
        RECT 72.365 39.630 72.645 40.630 ;
        RECT 74.675 37.655 74.955 40.630 ;
        RECT 76.925 39.630 77.205 40.630 ;
        RECT 78.205 39.630 78.485 40.630 ;
        RECT 79.485 39.630 79.765 40.630 ;
        RECT 80.765 39.630 81.045 40.630 ;
        RECT 82.045 39.630 82.325 40.630 ;
        RECT 70.115 37.325 74.955 37.655 ;
        RECT 66.280 36.420 66.860 36.750 ;
        RECT 64.640 35.730 64.930 36.230 ;
        RECT 65.275 35.730 65.555 36.230 ;
        RECT 64.640 32.990 64.930 33.490 ;
        RECT 65.675 32.990 65.955 33.490 ;
        RECT 66.280 31.745 66.610 36.420 ;
        RECT 67.835 34.755 68.115 36.230 ;
        RECT 70.115 35.730 70.395 37.325 ;
        RECT 72.395 34.755 72.675 36.230 ;
        RECT 74.675 35.730 74.955 37.325 ;
        RECT 84.355 38.480 84.635 40.630 ;
        RECT 86.605 39.630 86.885 40.630 ;
        RECT 87.885 39.630 88.165 40.630 ;
        RECT 89.165 39.630 89.445 40.630 ;
        RECT 89.830 39.630 90.120 40.630 ;
        RECT 84.355 38.150 89.195 38.480 ;
        RECT 76.955 34.755 77.235 36.230 ;
        RECT 78.235 35.730 78.515 36.230 ;
        RECT 79.515 35.730 79.795 36.230 ;
        RECT 80.795 35.730 81.075 36.230 ;
        RECT 82.075 34.755 82.355 36.230 ;
        RECT 84.355 35.730 84.635 38.150 ;
        RECT 86.635 34.755 86.915 36.230 ;
        RECT 88.915 35.730 89.195 38.150 ;
        RECT 92.700 36.750 93.030 47.530 ;
        RECT 94.080 44.475 94.370 45.475 ;
        RECT 94.755 44.475 95.035 45.475 ;
        RECT 97.035 44.475 97.315 45.475 ;
        RECT 99.315 44.475 99.595 45.475 ;
        RECT 99.760 43.955 100.660 44.285 ;
        RECT 100.070 42.790 100.350 43.955 ;
        RECT 99.625 42.460 100.795 42.790 ;
        RECT 99.625 41.780 100.795 42.110 ;
        RECT 100.070 41.195 100.350 41.780 ;
        RECT 99.760 40.865 100.660 41.195 ;
        RECT 94.080 40.175 94.370 40.675 ;
        RECT 94.755 40.175 95.035 40.675 ;
        RECT 97.035 40.175 97.315 40.675 ;
        RECT 99.315 40.175 99.595 40.675 ;
        RECT 101.595 40.175 101.875 45.475 ;
        RECT 103.875 44.475 104.155 45.475 ;
        RECT 103.875 40.175 104.155 40.675 ;
        RECT 106.155 40.175 106.435 45.475 ;
        RECT 108.435 44.475 108.715 45.475 ;
        RECT 108.435 40.175 108.715 40.675 ;
        RECT 110.715 40.175 110.995 45.475 ;
        RECT 112.995 44.475 113.275 45.475 ;
        RECT 115.275 44.475 115.555 45.475 ;
        RECT 117.555 44.475 117.835 45.475 ;
        RECT 118.220 44.475 118.510 45.475 ;
        RECT 112.995 40.175 113.275 40.675 ;
        RECT 115.275 40.175 115.555 40.675 ;
        RECT 117.555 40.175 117.835 40.675 ;
        RECT 118.220 40.175 118.510 40.675 ;
        RECT 92.450 36.420 93.030 36.750 ;
        RECT 91.195 34.755 91.475 36.230 ;
        RECT 67.635 34.385 68.315 34.755 ;
        RECT 72.195 34.385 72.875 34.755 ;
        RECT 76.755 34.385 77.435 34.755 ;
        RECT 79.070 34.405 80.240 34.735 ;
        RECT 68.955 32.990 69.235 33.490 ;
        RECT 72.235 32.990 72.515 33.490 ;
        RECT 79.515 32.990 79.795 34.405 ;
        RECT 81.875 34.385 82.555 34.755 ;
        RECT 86.435 34.385 87.115 34.755 ;
        RECT 90.995 34.385 91.675 34.755 ;
        RECT 86.795 32.990 87.075 33.490 ;
        RECT 90.075 32.990 90.355 33.490 ;
        RECT 80.605 32.470 81.825 32.800 ;
        RECT 80.715 31.960 81.715 32.470 ;
        RECT 65.505 31.145 66.610 31.745 ;
        RECT 65.505 29.045 66.610 29.645 ;
        RECT 64.640 27.300 64.930 27.800 ;
        RECT 65.675 27.300 65.955 27.800 ;
        RECT 64.640 24.560 64.930 25.060 ;
        RECT 65.275 24.560 65.555 25.060 ;
        RECT 66.280 24.370 66.610 29.045 ;
        RECT 80.715 28.320 81.715 28.830 ;
        RECT 80.605 27.990 81.825 28.320 ;
        RECT 68.955 27.300 69.235 27.800 ;
        RECT 72.235 27.300 72.515 27.800 ;
        RECT 67.635 26.035 68.315 26.405 ;
        RECT 72.195 26.035 72.875 26.405 ;
        RECT 76.755 26.035 77.435 26.405 ;
        RECT 79.515 26.385 79.795 27.800 ;
        RECT 86.795 27.300 87.075 27.800 ;
        RECT 90.075 27.300 90.355 27.800 ;
        RECT 79.070 26.055 80.240 26.385 ;
        RECT 81.875 26.035 82.555 26.405 ;
        RECT 86.435 26.035 87.115 26.405 ;
        RECT 90.995 26.035 91.675 26.405 ;
        RECT 67.835 24.560 68.115 26.035 ;
        RECT 66.280 24.040 66.860 24.370 ;
        RECT 60.435 23.135 61.605 23.465 ;
        RECT 55.440 22.310 56.610 22.640 ;
        RECT 55.440 14.150 55.720 22.310 ;
        RECT 55.920 16.405 56.210 16.905 ;
        RECT 56.595 16.405 56.875 16.905 ;
        RECT 57.375 16.405 57.655 16.905 ;
        RECT 58.155 16.405 58.435 16.905 ;
        RECT 60.435 16.405 60.715 23.135 ;
        RECT 62.715 16.405 62.995 16.905 ;
        RECT 63.495 16.405 63.775 16.905 ;
        RECT 64.275 16.405 64.555 16.905 ;
        RECT 64.940 16.405 65.230 16.905 ;
        RECT 60.125 15.885 61.025 16.215 ;
        RECT 60.435 15.095 60.715 15.885 ;
        RECT 60.435 14.765 61.605 15.095 ;
        RECT 57.720 14.170 58.890 14.500 ;
        RECT 58.600 13.260 58.890 14.170 ;
        RECT 58.600 12.930 59.500 13.260 ;
        RECT 55.920 11.740 56.210 12.740 ;
        RECT 56.595 11.740 56.875 12.740 ;
        RECT 57.375 11.740 57.655 12.740 ;
        RECT 58.155 11.740 58.435 12.740 ;
        RECT 60.435 11.740 60.715 14.435 ;
        RECT 66.280 13.260 66.610 24.040 ;
        RECT 70.115 23.465 70.395 25.060 ;
        RECT 72.395 24.560 72.675 26.035 ;
        RECT 74.675 23.465 74.955 25.060 ;
        RECT 76.955 24.560 77.235 26.035 ;
        RECT 78.235 24.560 78.515 25.060 ;
        RECT 79.515 24.560 79.795 25.060 ;
        RECT 80.795 24.560 81.075 25.060 ;
        RECT 82.075 24.560 82.355 26.035 ;
        RECT 70.115 23.135 74.955 23.465 ;
        RECT 69.130 20.160 69.420 21.160 ;
        RECT 69.805 20.160 70.085 21.160 ;
        RECT 71.085 20.160 71.365 21.160 ;
        RECT 72.365 20.160 72.645 21.160 ;
        RECT 74.675 20.160 74.955 23.135 ;
        RECT 84.355 22.640 84.635 25.060 ;
        RECT 86.635 24.560 86.915 26.035 ;
        RECT 88.915 22.640 89.195 25.060 ;
        RECT 91.195 24.560 91.475 26.035 ;
        RECT 92.700 24.370 93.030 36.420 ;
        RECT 93.755 35.730 94.035 36.230 ;
        RECT 94.380 35.730 94.670 36.230 ;
        RECT 93.355 32.990 93.635 33.490 ;
        RECT 94.380 32.990 94.670 33.490 ;
        RECT 120.560 30.165 121.160 55.070 ;
        RECT 124.400 43.960 124.690 44.960 ;
        RECT 125.075 43.960 125.355 44.960 ;
        RECT 125.505 43.960 125.785 44.960 ;
        RECT 125.935 43.960 126.215 44.960 ;
        RECT 126.365 42.450 126.645 45.460 ;
        RECT 126.795 43.960 127.075 44.960 ;
        RECT 127.225 42.450 127.505 45.460 ;
        RECT 127.655 43.960 127.935 44.960 ;
        RECT 128.085 43.960 128.365 44.960 ;
        RECT 128.515 43.960 128.795 44.960 ;
        RECT 129.180 43.960 129.470 44.960 ;
        RECT 132.225 42.450 132.555 46.795 ;
        RECT 135.060 43.960 135.350 44.960 ;
        RECT 135.735 43.960 136.015 44.960 ;
        RECT 136.165 43.960 136.445 44.960 ;
        RECT 136.595 43.960 136.875 44.960 ;
        RECT 137.025 42.450 137.305 45.460 ;
        RECT 137.455 43.960 137.735 44.960 ;
        RECT 137.885 42.450 138.165 45.460 ;
        RECT 138.315 43.960 138.595 44.960 ;
        RECT 125.085 42.120 125.855 42.450 ;
        RECT 126.365 42.120 130.740 42.450 ;
        RECT 132.225 42.120 133.395 42.450 ;
        RECT 135.745 42.120 136.515 42.450 ;
        RECT 137.025 42.120 138.165 42.450 ;
        RECT 124.400 40.110 124.690 41.110 ;
        RECT 125.075 40.110 125.355 41.110 ;
        RECT 125.505 40.110 125.785 41.110 ;
        RECT 125.935 40.110 126.215 41.110 ;
        RECT 126.365 40.110 126.645 42.120 ;
        RECT 126.795 40.110 127.075 41.110 ;
        RECT 127.225 40.110 127.505 42.120 ;
        RECT 127.655 40.110 127.935 41.110 ;
        RECT 128.085 40.110 128.365 41.110 ;
        RECT 128.515 40.110 128.795 41.110 ;
        RECT 129.180 40.110 129.470 41.110 ;
        RECT 130.410 39.005 130.740 42.120 ;
        RECT 135.060 40.110 135.350 41.110 ;
        RECT 135.735 40.110 136.015 41.110 ;
        RECT 136.165 40.110 136.445 41.110 ;
        RECT 136.595 40.110 136.875 41.110 ;
        RECT 137.025 40.110 137.305 42.120 ;
        RECT 137.455 40.110 137.735 41.110 ;
        RECT 137.885 40.110 138.165 42.120 ;
        RECT 138.745 42.450 139.025 45.460 ;
        RECT 139.175 43.960 139.455 44.960 ;
        RECT 139.605 42.450 139.885 45.460 ;
        RECT 140.035 43.960 140.315 44.960 ;
        RECT 140.465 42.450 140.745 45.460 ;
        RECT 140.895 43.960 141.175 44.960 ;
        RECT 141.325 42.450 141.605 45.460 ;
        RECT 141.755 43.960 142.035 44.960 ;
        RECT 142.185 42.450 142.465 45.460 ;
        RECT 142.615 43.960 142.895 44.960 ;
        RECT 143.045 43.960 143.325 44.960 ;
        RECT 143.475 43.960 143.755 44.960 ;
        RECT 144.140 43.960 144.430 44.960 ;
        RECT 138.745 42.120 143.700 42.450 ;
        RECT 138.315 40.110 138.595 41.110 ;
        RECT 138.745 40.110 139.025 42.120 ;
        RECT 139.175 40.110 139.455 41.110 ;
        RECT 139.605 40.110 139.885 42.120 ;
        RECT 140.035 40.110 140.315 41.110 ;
        RECT 140.465 40.110 140.745 42.120 ;
        RECT 140.895 40.110 141.175 41.110 ;
        RECT 141.325 40.110 141.605 42.120 ;
        RECT 141.755 40.110 142.035 41.110 ;
        RECT 142.185 40.110 142.465 42.120 ;
        RECT 142.615 40.110 142.895 41.110 ;
        RECT 143.045 40.110 143.325 41.110 ;
        RECT 143.475 40.110 143.755 41.110 ;
        RECT 144.140 40.110 144.430 41.110 ;
        RECT 122.365 38.675 130.740 39.005 ;
        RECT 122.365 34.780 122.695 38.675 ;
        RECT 93.355 27.300 93.635 27.800 ;
        RECT 94.380 27.300 94.670 27.800 ;
        RECT 123.495 25.410 123.825 38.435 ;
        RECT 129.125 38.085 130.295 38.415 ;
        RECT 124.125 37.305 125.295 37.635 ;
        RECT 124.125 30.975 124.405 37.305 ;
        RECT 126.515 37.285 127.195 37.655 ;
        RECT 124.750 36.115 125.040 36.965 ;
        RECT 125.425 36.115 125.705 36.965 ;
        RECT 125.855 36.115 126.135 36.965 ;
        RECT 126.285 36.115 126.565 36.965 ;
        RECT 126.715 35.130 126.995 37.115 ;
        RECT 127.145 36.115 127.425 36.965 ;
        RECT 127.575 35.130 127.855 37.115 ;
        RECT 128.005 36.115 128.285 36.965 ;
        RECT 128.435 36.115 128.715 36.965 ;
        RECT 128.865 36.115 129.145 36.965 ;
        RECT 129.515 36.115 129.820 36.965 ;
        RECT 129.965 35.130 130.295 38.085 ;
        RECT 135.060 36.140 135.350 37.140 ;
        RECT 135.735 36.140 136.015 37.140 ;
        RECT 136.165 36.140 136.445 37.140 ;
        RECT 136.595 36.140 136.875 37.140 ;
        RECT 137.025 35.130 137.305 37.140 ;
        RECT 137.455 36.140 137.735 37.140 ;
        RECT 137.885 35.130 138.165 37.140 ;
        RECT 138.315 36.140 138.595 37.140 ;
        RECT 125.505 34.800 126.365 35.130 ;
        RECT 126.715 34.800 130.295 35.130 ;
        RECT 135.745 34.800 136.515 35.130 ;
        RECT 137.025 34.800 138.165 35.130 ;
        RECT 124.750 32.890 125.040 33.740 ;
        RECT 125.425 32.890 125.705 33.740 ;
        RECT 125.855 32.890 126.135 33.740 ;
        RECT 126.285 32.635 126.565 33.815 ;
        RECT 126.715 32.815 126.995 34.800 ;
        RECT 127.145 32.635 127.425 33.815 ;
        RECT 127.575 32.815 127.855 34.800 ;
        RECT 128.005 32.635 128.285 33.815 ;
        RECT 128.435 32.890 128.715 33.740 ;
        RECT 128.865 32.890 129.145 33.740 ;
        RECT 129.515 32.890 129.820 33.740 ;
        RECT 126.285 32.345 128.285 32.635 ;
        RECT 124.750 31.315 125.040 32.165 ;
        RECT 125.425 31.315 125.705 32.165 ;
        RECT 125.855 31.315 126.135 32.165 ;
        RECT 126.285 31.315 126.565 32.165 ;
        RECT 126.715 31.165 126.995 32.345 ;
        RECT 127.145 31.315 127.425 32.165 ;
        RECT 127.575 31.165 127.855 32.345 ;
        RECT 135.060 32.290 135.350 33.290 ;
        RECT 135.735 32.290 136.015 33.290 ;
        RECT 136.165 32.290 136.445 33.290 ;
        RECT 136.595 32.290 136.875 33.290 ;
        RECT 128.005 31.315 128.285 32.165 ;
        RECT 128.435 31.315 128.715 32.165 ;
        RECT 128.865 31.315 129.145 32.165 ;
        RECT 129.515 31.315 129.820 32.165 ;
        RECT 137.025 31.790 137.305 34.800 ;
        RECT 137.455 32.290 137.735 33.290 ;
        RECT 137.885 31.790 138.165 34.800 ;
        RECT 138.745 35.130 139.025 37.140 ;
        RECT 139.175 36.140 139.455 37.140 ;
        RECT 139.605 35.130 139.885 37.140 ;
        RECT 140.035 36.140 140.315 37.140 ;
        RECT 140.465 35.130 140.745 37.140 ;
        RECT 140.895 36.140 141.175 37.140 ;
        RECT 141.325 35.130 141.605 37.140 ;
        RECT 141.755 36.140 142.035 37.140 ;
        RECT 142.185 35.130 142.465 37.140 ;
        RECT 142.615 36.140 142.895 37.140 ;
        RECT 143.045 36.140 143.325 37.140 ;
        RECT 143.475 36.140 143.755 37.140 ;
        RECT 144.140 36.140 144.430 37.140 ;
        RECT 138.745 34.800 143.700 35.130 ;
        RECT 138.315 32.290 138.595 33.290 ;
        RECT 138.745 31.790 139.025 34.800 ;
        RECT 139.175 32.290 139.455 33.290 ;
        RECT 139.605 31.790 139.885 34.800 ;
        RECT 140.035 32.290 140.315 33.290 ;
        RECT 140.465 31.790 140.745 34.800 ;
        RECT 140.895 32.290 141.175 33.290 ;
        RECT 141.325 31.790 141.605 34.800 ;
        RECT 141.755 32.290 142.035 33.290 ;
        RECT 142.185 31.790 142.465 34.800 ;
        RECT 142.615 32.290 142.895 33.290 ;
        RECT 143.045 32.290 143.325 33.290 ;
        RECT 143.475 32.290 143.755 33.290 ;
        RECT 144.140 32.290 144.430 33.290 ;
        RECT 124.125 30.645 125.295 30.975 ;
        RECT 126.560 30.645 128.010 30.975 ;
        RECT 124.125 30.565 124.405 30.645 ;
        RECT 124.125 29.915 124.405 29.995 ;
        RECT 124.125 29.585 125.295 29.915 ;
        RECT 126.560 29.585 128.010 29.915 ;
        RECT 93.755 24.560 94.035 25.060 ;
        RECT 94.380 24.560 94.670 25.060 ;
        RECT 92.450 24.040 93.030 24.370 ;
        RECT 84.355 22.310 89.195 22.640 ;
        RECT 76.925 20.160 77.205 21.160 ;
        RECT 78.205 20.160 78.485 21.160 ;
        RECT 79.485 20.160 79.765 21.160 ;
        RECT 80.765 20.160 81.045 21.160 ;
        RECT 82.045 20.160 82.325 21.160 ;
        RECT 84.355 20.160 84.635 22.310 ;
        RECT 86.605 20.160 86.885 21.160 ;
        RECT 87.885 20.160 88.165 21.160 ;
        RECT 89.165 20.160 89.445 21.160 ;
        RECT 89.830 20.160 90.120 21.160 ;
        RECT 75.860 19.640 76.760 19.970 ;
        RECT 73.120 18.680 74.290 19.010 ;
        RECT 73.120 17.425 73.400 18.680 ;
        RECT 76.170 18.330 76.450 19.640 ;
        RECT 75.280 18.000 76.450 18.330 ;
        RECT 72.810 17.095 73.710 17.425 ;
        RECT 69.130 16.405 69.420 16.905 ;
        RECT 69.805 16.405 70.085 16.905 ;
        RECT 71.085 16.405 71.365 16.905 ;
        RECT 72.365 16.405 72.645 16.905 ;
        RECT 76.925 16.405 77.205 16.905 ;
        RECT 78.205 16.405 78.485 16.905 ;
        RECT 79.485 16.405 79.765 16.905 ;
        RECT 80.765 16.405 81.045 16.905 ;
        RECT 82.045 16.405 82.325 16.905 ;
        RECT 72.675 15.885 73.575 16.215 ;
        RECT 84.325 16.210 84.605 16.905 ;
        RECT 86.605 16.405 86.885 16.905 ;
        RECT 87.885 16.405 88.165 16.905 ;
        RECT 89.165 16.405 89.445 16.905 ;
        RECT 89.830 16.405 90.120 16.905 ;
        RECT 66.280 12.930 67.180 13.260 ;
        RECT 62.715 11.740 62.995 12.740 ;
        RECT 63.495 11.740 63.775 12.740 ;
        RECT 64.275 11.740 64.555 12.740 ;
        RECT 65.055 11.740 65.335 12.740 ;
        RECT 65.835 10.585 66.115 12.740 ;
        RECT 68.115 11.740 68.395 14.435 ;
        RECT 70.395 10.585 70.675 12.740 ;
        RECT 72.675 11.740 72.955 15.885 ;
        RECT 84.015 15.880 84.915 16.210 ;
        RECT 84.325 15.095 84.605 15.880 ;
        RECT 83.435 14.765 84.605 15.095 ;
        RECT 74.955 10.585 75.235 12.740 ;
        RECT 77.235 11.740 77.515 14.435 ;
        RECT 79.515 10.585 79.795 12.740 ;
        RECT 81.795 11.740 82.075 14.435 ;
        RECT 84.325 14.415 84.605 14.765 ;
        RECT 83.880 14.085 85.050 14.415 ;
        RECT 84.075 10.585 84.355 12.740 ;
        RECT 86.355 11.740 86.635 14.435 ;
        RECT 88.635 10.585 88.915 12.740 ;
        RECT 90.915 11.740 91.195 14.435 ;
        RECT 92.700 13.260 93.030 24.040 ;
        RECT 124.125 23.255 124.405 29.585 ;
        RECT 124.750 28.395 125.040 29.245 ;
        RECT 125.425 28.395 125.705 29.245 ;
        RECT 125.855 28.395 126.135 29.245 ;
        RECT 126.285 28.395 126.565 29.245 ;
        RECT 126.715 28.215 126.995 29.395 ;
        RECT 127.145 28.395 127.425 29.245 ;
        RECT 127.575 28.215 127.855 29.395 ;
        RECT 128.005 28.395 128.285 29.245 ;
        RECT 128.435 28.395 128.715 29.245 ;
        RECT 128.865 28.395 129.145 29.245 ;
        RECT 129.515 28.395 129.820 29.245 ;
        RECT 126.285 27.925 128.285 28.215 ;
        RECT 124.750 26.820 125.040 27.670 ;
        RECT 125.425 26.820 125.705 27.670 ;
        RECT 125.855 26.820 126.135 27.670 ;
        RECT 126.285 26.745 126.565 27.925 ;
        RECT 126.715 25.760 126.995 27.745 ;
        RECT 127.145 26.745 127.425 27.925 ;
        RECT 127.575 25.760 127.855 27.745 ;
        RECT 128.005 26.745 128.285 27.925 ;
        RECT 129.965 27.690 130.295 30.995 ;
        RECT 135.060 29.200 135.350 30.200 ;
        RECT 135.735 29.200 136.015 30.200 ;
        RECT 136.165 29.200 136.445 30.200 ;
        RECT 136.595 29.200 136.875 30.200 ;
        RECT 137.025 27.690 137.305 30.700 ;
        RECT 137.455 29.200 137.735 30.200 ;
        RECT 137.885 27.690 138.165 30.700 ;
        RECT 138.315 29.200 138.595 30.200 ;
        RECT 128.435 26.820 128.715 27.670 ;
        RECT 128.865 26.820 129.145 27.670 ;
        RECT 129.515 26.820 129.820 27.670 ;
        RECT 129.965 27.360 131.970 27.690 ;
        RECT 135.745 27.360 136.515 27.690 ;
        RECT 137.025 27.360 138.165 27.690 ;
        RECT 129.965 25.760 130.295 27.360 ;
        RECT 125.505 25.430 126.365 25.760 ;
        RECT 126.715 25.430 130.295 25.760 ;
        RECT 124.750 23.595 125.040 24.445 ;
        RECT 125.425 23.595 125.705 24.445 ;
        RECT 125.855 23.595 126.135 24.445 ;
        RECT 126.285 23.595 126.565 24.445 ;
        RECT 126.715 23.445 126.995 25.430 ;
        RECT 127.145 23.595 127.425 24.445 ;
        RECT 127.575 23.445 127.855 25.430 ;
        RECT 135.060 25.350 135.350 26.350 ;
        RECT 135.735 25.350 136.015 26.350 ;
        RECT 136.165 25.350 136.445 26.350 ;
        RECT 136.595 25.350 136.875 26.350 ;
        RECT 137.025 25.350 137.305 27.360 ;
        RECT 137.455 25.350 137.735 26.350 ;
        RECT 137.885 25.350 138.165 27.360 ;
        RECT 138.745 27.690 139.025 30.700 ;
        RECT 139.175 29.200 139.455 30.200 ;
        RECT 139.605 27.690 139.885 30.700 ;
        RECT 140.035 29.200 140.315 30.200 ;
        RECT 140.465 27.690 140.745 30.700 ;
        RECT 140.895 29.200 141.175 30.200 ;
        RECT 141.325 27.690 141.605 30.700 ;
        RECT 141.755 29.200 142.035 30.200 ;
        RECT 142.185 27.690 142.465 30.700 ;
        RECT 142.615 29.200 142.895 30.200 ;
        RECT 143.045 29.200 143.325 30.200 ;
        RECT 143.475 29.200 143.755 30.200 ;
        RECT 144.140 29.200 144.430 30.200 ;
        RECT 138.745 27.360 143.700 27.690 ;
        RECT 138.315 25.350 138.595 26.350 ;
        RECT 138.745 25.350 139.025 27.360 ;
        RECT 139.175 25.350 139.455 26.350 ;
        RECT 139.605 25.350 139.885 27.360 ;
        RECT 140.035 25.350 140.315 26.350 ;
        RECT 140.465 25.350 140.745 27.360 ;
        RECT 140.895 25.350 141.175 26.350 ;
        RECT 141.325 25.350 141.605 27.360 ;
        RECT 141.755 25.350 142.035 26.350 ;
        RECT 142.185 25.350 142.465 27.360 ;
        RECT 142.615 25.350 142.895 26.350 ;
        RECT 143.045 25.350 143.325 26.350 ;
        RECT 143.475 25.350 143.755 26.350 ;
        RECT 144.140 25.350 144.430 26.350 ;
        RECT 128.005 23.595 128.285 24.445 ;
        RECT 128.435 23.595 128.715 24.445 ;
        RECT 128.865 23.595 129.145 24.445 ;
        RECT 129.515 23.595 129.820 24.445 ;
        RECT 187.345 23.610 187.675 74.960 ;
        RECT 188.175 38.515 188.505 74.375 ;
        RECT 189.005 56.170 189.605 69.045 ;
        RECT 194.205 68.715 194.805 93.530 ;
        RECT 202.970 85.480 203.570 108.665 ;
        RECT 190.690 41.985 191.770 42.585 ;
        RECT 186.505 23.280 187.675 23.610 ;
        RECT 124.125 22.925 125.295 23.255 ;
        RECT 126.515 22.905 127.195 23.275 ;
        RECT 94.080 20.115 94.370 20.615 ;
        RECT 94.755 20.115 95.035 20.615 ;
        RECT 97.035 20.115 97.315 20.615 ;
        RECT 99.315 20.115 99.595 20.615 ;
        RECT 99.760 19.595 100.660 19.925 ;
        RECT 100.070 19.010 100.350 19.595 ;
        RECT 99.625 18.680 100.795 19.010 ;
        RECT 99.625 18.000 100.795 18.330 ;
        RECT 100.070 16.835 100.350 18.000 ;
        RECT 99.760 16.505 100.660 16.835 ;
        RECT 94.080 15.315 94.370 16.315 ;
        RECT 94.755 15.315 95.035 16.315 ;
        RECT 97.035 15.315 97.315 16.315 ;
        RECT 99.315 15.315 99.595 16.315 ;
        RECT 101.595 15.315 101.875 20.615 ;
        RECT 103.875 20.115 104.155 20.615 ;
        RECT 103.875 15.315 104.155 16.315 ;
        RECT 106.155 15.315 106.435 20.615 ;
        RECT 108.435 20.115 108.715 20.615 ;
        RECT 108.435 15.315 108.715 16.315 ;
        RECT 110.715 15.315 110.995 20.615 ;
        RECT 112.995 20.115 113.275 20.615 ;
        RECT 115.275 20.115 115.555 20.615 ;
        RECT 117.555 20.115 117.835 20.615 ;
        RECT 118.220 20.115 118.510 20.615 ;
        RECT 135.060 20.180 135.350 21.180 ;
        RECT 135.735 20.180 136.015 21.180 ;
        RECT 136.165 20.180 136.445 21.180 ;
        RECT 136.595 20.180 136.875 21.180 ;
        RECT 137.025 18.670 137.305 21.680 ;
        RECT 137.455 20.180 137.735 21.180 ;
        RECT 137.885 18.670 138.165 21.680 ;
        RECT 138.315 20.180 138.595 21.180 ;
        RECT 135.745 18.340 136.515 18.670 ;
        RECT 137.025 18.340 138.165 18.670 ;
        RECT 135.060 16.330 135.350 17.330 ;
        RECT 135.735 16.330 136.015 17.330 ;
        RECT 136.165 16.330 136.445 17.330 ;
        RECT 136.595 16.330 136.875 17.330 ;
        RECT 137.025 16.330 137.305 18.340 ;
        RECT 137.455 16.330 137.735 17.330 ;
        RECT 137.885 16.330 138.165 18.340 ;
        RECT 138.745 18.670 139.025 21.680 ;
        RECT 139.175 20.180 139.455 21.180 ;
        RECT 139.605 18.670 139.885 21.680 ;
        RECT 140.035 20.180 140.315 21.180 ;
        RECT 140.465 18.670 140.745 21.680 ;
        RECT 140.895 20.180 141.175 21.180 ;
        RECT 141.325 18.670 141.605 21.680 ;
        RECT 141.755 20.180 142.035 21.180 ;
        RECT 142.185 18.670 142.465 21.680 ;
        RECT 142.615 20.180 142.895 21.180 ;
        RECT 143.045 20.180 143.325 21.180 ;
        RECT 143.475 20.180 143.755 21.180 ;
        RECT 144.140 20.180 144.430 21.180 ;
        RECT 138.745 18.340 143.700 18.670 ;
        RECT 138.315 16.330 138.595 17.330 ;
        RECT 138.745 16.330 139.025 18.340 ;
        RECT 139.175 16.330 139.455 17.330 ;
        RECT 139.605 16.330 139.885 18.340 ;
        RECT 140.035 16.330 140.315 17.330 ;
        RECT 140.465 16.330 140.745 18.340 ;
        RECT 140.895 16.330 141.175 17.330 ;
        RECT 141.325 16.330 141.605 18.340 ;
        RECT 141.755 16.330 142.035 17.330 ;
        RECT 142.185 16.330 142.465 18.340 ;
        RECT 142.615 16.330 142.895 17.330 ;
        RECT 143.045 16.330 143.325 17.330 ;
        RECT 143.475 16.330 143.755 17.330 ;
        RECT 144.140 16.330 144.430 17.330 ;
        RECT 112.995 15.315 113.275 16.315 ;
        RECT 115.275 15.315 115.555 16.315 ;
        RECT 117.555 15.315 117.835 16.315 ;
        RECT 118.220 15.315 118.510 16.315 ;
        RECT 92.130 12.930 93.030 13.260 ;
        RECT 93.195 10.585 93.475 12.740 ;
        RECT 93.975 11.740 94.255 12.740 ;
        RECT 94.755 11.740 95.035 12.740 ;
        RECT 95.420 11.740 95.710 12.740 ;
        RECT 65.835 10.255 93.475 10.585 ;
        RECT 55.920 8.150 56.210 9.150 ;
        RECT 65.835 8.150 66.115 9.150 ;
        RECT 68.115 8.150 68.395 9.150 ;
        RECT 70.395 8.150 70.675 9.150 ;
        RECT 72.675 8.150 72.955 9.150 ;
        RECT 74.955 8.150 75.235 9.150 ;
        RECT 77.235 8.150 77.515 9.150 ;
        RECT 79.515 8.150 79.795 10.255 ;
        RECT 81.795 8.150 82.075 9.150 ;
        RECT 84.075 8.150 84.355 9.150 ;
        RECT 86.355 8.150 86.635 9.150 ;
        RECT 88.635 8.150 88.915 9.150 ;
        RECT 90.915 8.150 91.195 9.150 ;
        RECT 93.195 8.150 93.475 9.150 ;
        RECT 95.420 8.150 95.710 9.150 ;
        RECT 79.205 7.630 80.105 7.960 ;
        RECT 79.490 7.430 79.820 7.630 ;
        RECT 78.650 7.100 79.820 7.430 ;
        RECT 191.170 -1.305 191.770 41.985 ;
        RECT 34.425 -1.905 191.770 -1.305 ;
        RECT 192.270 -2.405 192.870 35.265 ;
        RECT 199.550 27.225 200.150 64.000 ;
        RECT 200.650 18.205 201.250 41.920 ;
        RECT 33.325 -3.005 192.870 -2.405 ;
      LAYER via2 ;
        RECT -4.050 108.825 -3.770 109.105 ;
        RECT -3.650 108.825 -3.370 109.105 ;
        RECT -3.250 108.825 -2.970 109.105 ;
        RECT 202.090 108.825 202.370 109.105 ;
        RECT 202.490 108.825 202.770 109.105 ;
        RECT 202.890 108.825 203.170 109.105 ;
        RECT 203.290 108.825 203.570 109.105 ;
        RECT -4.855 94.830 -4.575 95.110 ;
        RECT -4.855 94.430 -4.575 94.710 ;
        RECT -4.855 94.030 -4.575 94.310 ;
        RECT -4.855 79.220 -4.575 79.500 ;
        RECT -4.855 78.820 -4.575 79.100 ;
        RECT -4.855 78.420 -4.575 78.700 ;
        RECT -2.390 107.725 -2.110 108.005 ;
        RECT -1.990 107.725 -1.710 108.005 ;
        RECT -3.195 98.505 -2.915 98.785 ;
        RECT -3.195 98.105 -2.915 98.385 ;
        RECT -3.195 97.705 -2.915 97.985 ;
        RECT -2.230 75.105 -1.950 75.385 ;
        RECT -2.230 74.705 -1.950 74.985 ;
        RECT -1.130 93.025 -0.850 93.305 ;
        RECT -1.130 92.625 -0.850 92.905 ;
        RECT -1.130 92.225 -0.850 92.505 ;
        RECT -1.130 91.825 -0.850 92.105 ;
        RECT -3.195 72.180 -2.915 72.460 ;
        RECT -3.195 71.780 -2.915 72.060 ;
        RECT -3.195 71.380 -2.915 71.660 ;
        RECT 168.765 93.025 169.045 93.305 ;
        RECT 168.765 92.625 169.045 92.905 ;
        RECT 168.765 92.225 169.045 92.505 ;
        RECT 168.765 91.825 169.045 92.105 ;
        RECT 141.660 78.420 141.940 78.700 ;
        RECT 142.060 78.420 142.340 78.700 ;
        RECT 142.460 78.420 142.740 78.700 ;
        RECT 137.115 76.635 137.395 76.915 ;
        RECT 137.745 76.635 138.025 76.915 ;
        RECT 138.175 76.635 138.455 76.915 ;
        RECT 138.605 76.635 138.885 76.915 ;
        RECT 139.035 76.635 139.315 76.915 ;
        RECT 139.465 76.635 139.745 76.915 ;
        RECT 139.895 76.635 140.175 76.915 ;
        RECT 140.325 76.635 140.605 76.915 ;
        RECT 140.755 76.635 141.035 76.915 ;
        RECT 141.185 76.635 141.465 76.915 ;
        RECT 142.045 76.635 142.325 76.915 ;
        RECT 142.905 76.635 143.185 76.915 ;
        RECT 143.335 76.635 143.615 76.915 ;
        RECT 143.765 76.635 144.045 76.915 ;
        RECT 144.195 76.635 144.475 76.915 ;
        RECT 144.625 76.635 144.905 76.915 ;
        RECT 145.055 76.635 145.335 76.915 ;
        RECT 145.485 76.635 145.765 76.915 ;
        RECT 145.915 76.635 146.195 76.915 ;
        RECT 146.345 76.635 146.625 76.915 ;
        RECT 146.975 76.635 147.255 76.915 ;
        RECT 168.765 76.465 169.045 76.745 ;
        RECT 42.715 75.390 42.995 75.670 ;
        RECT 43.345 75.390 43.625 75.670 ;
        RECT 45.625 75.390 45.905 75.670 ;
        RECT 50.185 75.390 50.465 75.670 ;
        RECT 54.745 75.390 55.025 75.670 ;
        RECT 59.305 75.390 59.585 75.670 ;
        RECT 63.865 75.390 64.145 75.670 ;
        RECT 68.425 75.390 68.705 75.670 ;
        RECT 72.985 75.390 73.265 75.670 ;
        RECT 77.545 75.390 77.825 75.670 ;
        RECT 82.105 75.390 82.385 75.670 ;
        RECT 41.190 74.705 41.470 74.985 ;
        RECT 41.590 74.705 41.870 74.985 ;
        RECT 41.990 74.705 42.270 74.985 ;
        RECT 42.715 74.020 42.995 74.300 ;
        RECT 43.345 74.020 43.625 74.300 ;
        RECT 45.625 74.020 45.905 74.300 ;
        RECT 50.185 74.020 50.465 74.300 ;
        RECT 54.745 74.020 55.025 74.300 ;
        RECT 59.305 74.020 59.585 74.300 ;
        RECT 63.865 74.020 64.145 74.300 ;
        RECT 68.425 74.020 68.705 74.300 ;
        RECT 72.985 74.020 73.265 74.300 ;
        RECT 77.545 74.020 77.825 74.300 ;
        RECT 82.105 74.020 82.385 74.300 ;
        RECT 86.665 75.390 86.945 75.670 ;
        RECT 86.665 74.020 86.945 74.300 ;
        RECT 91.225 75.390 91.505 75.670 ;
        RECT 91.225 74.020 91.505 74.300 ;
        RECT 95.785 75.390 96.065 75.670 ;
        RECT 95.785 74.020 96.065 74.300 ;
        RECT 100.345 75.390 100.625 75.670 ;
        RECT 100.345 74.020 100.625 74.300 ;
        RECT 104.905 75.390 105.185 75.670 ;
        RECT 104.905 74.020 105.185 74.300 ;
        RECT 109.465 75.390 109.745 75.670 ;
        RECT 109.465 74.020 109.745 74.300 ;
        RECT 114.025 75.390 114.305 75.670 ;
        RECT 114.025 74.020 114.305 74.300 ;
        RECT 118.585 75.390 118.865 75.670 ;
        RECT 120.865 75.390 121.145 75.670 ;
        RECT 123.145 75.390 123.425 75.670 ;
        RECT 125.425 75.390 125.705 75.670 ;
        RECT 127.705 75.390 127.985 75.670 ;
        RECT 129.985 75.390 130.265 75.670 ;
        RECT 130.615 75.390 130.895 75.670 ;
        RECT 150.170 75.800 150.450 76.080 ;
        RECT 150.570 75.800 150.850 76.080 ;
        RECT 150.970 75.800 151.250 76.080 ;
        RECT 151.370 75.800 151.650 76.080 ;
        RECT 151.770 75.800 152.050 76.080 ;
        RECT 168.765 76.065 169.045 76.345 ;
        RECT 194.365 93.025 194.645 93.305 ;
        RECT 194.365 92.625 194.645 92.905 ;
        RECT 194.365 92.225 194.645 92.505 ;
        RECT 194.365 91.825 194.645 92.105 ;
        RECT 168.765 75.665 169.045 75.945 ;
        RECT 185.955 75.800 186.235 76.080 ;
        RECT 186.355 75.800 186.635 76.080 ;
        RECT 186.755 75.800 187.035 76.080 ;
        RECT 136.165 74.985 136.445 75.265 ;
        RECT 136.565 74.985 136.845 75.265 ;
        RECT 136.965 74.985 137.245 75.265 ;
        RECT 118.585 74.020 118.865 74.300 ;
        RECT 120.865 74.020 121.145 74.300 ;
        RECT 123.145 74.020 123.425 74.300 ;
        RECT 93.170 71.380 93.450 71.660 ;
        RECT 93.570 71.380 93.850 71.660 ;
        RECT 93.970 71.380 94.250 71.660 ;
        RECT -1.130 69.540 -0.850 69.820 ;
        RECT -1.130 69.140 -0.850 69.420 ;
        RECT -1.130 68.740 -0.850 69.020 ;
        RECT 0.605 68.740 0.885 69.020 ;
        RECT 1.005 68.740 1.285 69.020 ;
        RECT 1.405 68.740 1.685 69.020 ;
        RECT -4.025 67.200 -3.745 67.480 ;
        RECT -4.025 66.800 -3.745 67.080 ;
        RECT -4.025 66.400 -3.745 66.680 ;
        RECT 90.925 68.740 91.205 69.020 ;
        RECT 91.325 68.740 91.605 69.020 ;
        RECT 91.725 68.740 92.005 69.020 ;
        RECT 92.125 68.740 92.405 69.020 ;
        RECT 92.525 68.740 92.805 69.020 ;
        RECT 92.925 68.740 93.205 69.020 ;
        RECT 93.325 68.740 93.605 69.020 ;
        RECT 93.725 68.740 94.005 69.020 ;
        RECT 94.125 68.740 94.405 69.020 ;
        RECT 94.525 68.740 94.805 69.020 ;
        RECT 94.925 68.740 95.205 69.020 ;
        RECT 95.325 68.740 95.605 69.020 ;
        RECT 95.725 68.740 96.005 69.020 ;
        RECT 96.125 68.740 96.405 69.020 ;
        RECT 39.670 67.810 39.950 68.090 ;
        RECT 40.070 67.810 40.350 68.090 ;
        RECT 40.470 67.810 40.750 68.090 ;
        RECT 33.525 63.605 33.805 63.885 ;
        RECT 33.525 63.205 33.805 63.485 ;
        RECT 34.195 63.605 34.475 63.885 ;
        RECT 34.195 63.205 34.475 63.485 ;
        RECT 34.625 63.605 34.905 63.885 ;
        RECT 34.625 63.205 34.905 63.485 ;
        RECT 35.055 63.605 35.335 63.885 ;
        RECT 35.055 63.205 35.335 63.485 ;
        RECT 35.915 63.605 36.195 63.885 ;
        RECT 35.915 63.205 36.195 63.485 ;
        RECT 36.775 63.605 37.055 63.885 ;
        RECT 36.775 63.205 37.055 63.485 ;
        RECT 37.205 63.605 37.485 63.885 ;
        RECT 37.205 63.205 37.485 63.485 ;
        RECT 37.635 63.605 37.915 63.885 ;
        RECT 37.635 63.205 37.915 63.485 ;
        RECT 38.305 63.605 38.585 63.885 ;
        RECT 38.305 63.205 38.585 63.485 ;
        RECT 34.250 61.230 34.530 61.510 ;
        RECT 34.650 61.230 34.930 61.510 ;
        RECT 90.265 66.400 90.545 66.680 ;
        RECT 90.665 66.400 90.945 66.680 ;
        RECT 96.815 67.810 97.095 68.090 ;
        RECT 97.215 67.810 97.495 68.090 ;
        RECT 106.425 65.310 106.705 65.590 ;
        RECT 106.825 65.310 107.105 65.590 ;
        RECT 107.225 65.310 107.505 65.590 ;
        RECT 42.675 63.555 42.955 63.835 ;
        RECT 43.345 63.555 43.625 63.835 ;
        RECT 45.625 63.555 45.905 63.835 ;
        RECT 47.905 63.555 48.185 63.835 ;
        RECT 52.465 63.555 52.745 63.835 ;
        RECT 57.025 63.555 57.305 63.835 ;
        RECT 61.585 63.555 61.865 63.835 ;
        RECT 66.145 63.555 66.425 63.835 ;
        RECT 70.705 63.555 70.985 63.835 ;
        RECT 42.675 62.185 42.955 62.465 ;
        RECT 43.345 62.185 43.625 62.465 ;
        RECT 45.625 62.185 45.905 62.465 ;
        RECT 47.905 62.185 48.185 62.465 ;
        RECT 37.085 61.230 37.365 61.510 ;
        RECT 37.485 61.230 37.765 61.510 ;
        RECT 52.465 62.185 52.745 62.465 ;
        RECT 57.025 62.185 57.305 62.465 ;
        RECT 61.585 62.185 61.865 62.465 ;
        RECT 66.145 62.185 66.425 62.465 ;
        RECT 70.705 62.185 70.985 62.465 ;
        RECT 33.525 59.755 33.805 60.035 ;
        RECT 33.525 59.355 33.805 59.635 ;
        RECT 34.195 59.755 34.475 60.035 ;
        RECT 34.195 59.355 34.475 59.635 ;
        RECT 34.625 59.755 34.905 60.035 ;
        RECT 34.625 59.355 34.905 59.635 ;
        RECT 35.055 59.755 35.335 60.035 ;
        RECT 35.055 59.355 35.335 59.635 ;
        RECT 35.915 59.755 36.195 60.035 ;
        RECT 35.915 59.355 36.195 59.635 ;
        RECT 42.675 60.815 42.955 61.095 ;
        RECT 43.345 60.815 43.625 61.095 ;
        RECT 45.625 60.815 45.905 61.095 ;
        RECT 47.905 60.815 48.185 61.095 ;
        RECT 52.465 60.815 52.745 61.095 ;
        RECT 57.025 60.815 57.305 61.095 ;
        RECT 61.585 60.815 61.865 61.095 ;
        RECT 66.145 60.815 66.425 61.095 ;
        RECT 70.705 60.815 70.985 61.095 ;
        RECT 75.265 63.555 75.545 63.835 ;
        RECT 75.265 62.185 75.545 62.465 ;
        RECT 75.265 60.815 75.545 61.095 ;
        RECT 79.825 63.555 80.105 63.835 ;
        RECT 79.825 62.185 80.105 62.465 ;
        RECT 79.825 60.815 80.105 61.095 ;
        RECT 84.385 63.555 84.665 63.835 ;
        RECT 84.385 62.185 84.665 62.465 ;
        RECT 84.385 60.815 84.665 61.095 ;
        RECT 88.945 63.555 89.225 63.835 ;
        RECT 88.945 62.185 89.225 62.465 ;
        RECT 88.945 60.815 89.225 61.095 ;
        RECT 93.505 63.555 93.785 63.835 ;
        RECT 93.505 62.185 93.785 62.465 ;
        RECT 93.505 60.815 93.785 61.095 ;
        RECT 98.065 63.555 98.345 63.835 ;
        RECT 98.065 62.185 98.345 62.465 ;
        RECT 98.065 60.815 98.345 61.095 ;
        RECT 102.625 63.555 102.905 63.835 ;
        RECT 102.625 62.185 102.905 62.465 ;
        RECT 102.625 60.815 102.905 61.095 ;
        RECT 107.185 63.555 107.465 63.835 ;
        RECT 127.705 74.020 127.985 74.300 ;
        RECT 129.985 74.020 130.265 74.300 ;
        RECT 130.615 74.020 130.895 74.300 ;
        RECT 125.470 72.180 125.750 72.460 ;
        RECT 125.870 72.180 126.150 72.460 ;
        RECT 126.270 72.180 126.550 72.460 ;
        RECT 127.370 71.380 127.650 71.660 ;
        RECT 127.770 71.380 128.050 71.660 ;
        RECT 128.170 71.380 128.450 71.660 ;
        RECT 137.770 74.070 138.050 74.350 ;
        RECT 138.170 74.070 138.450 74.350 ;
        RECT 138.605 72.600 138.885 72.880 ;
        RECT 138.605 72.200 138.885 72.480 ;
        RECT 139.465 72.600 139.745 72.880 ;
        RECT 139.465 72.200 139.745 72.480 ;
        RECT 140.325 72.600 140.605 72.880 ;
        RECT 140.325 72.200 140.605 72.480 ;
        RECT 143.855 72.600 144.135 72.880 ;
        RECT 143.855 72.200 144.135 72.480 ;
        RECT 143.140 71.465 143.420 71.745 ;
        RECT 143.540 71.465 143.820 71.745 ;
        RECT 144.715 72.600 144.995 72.880 ;
        RECT 144.715 72.200 144.995 72.480 ;
        RECT 145.920 74.985 146.200 75.265 ;
        RECT 146.320 74.985 146.600 75.265 ;
        RECT 147.945 74.070 148.225 74.350 ;
        RECT 145.575 72.580 145.855 72.860 ;
        RECT 145.575 72.180 145.855 72.460 ;
        RECT 147.945 73.670 148.225 73.950 ;
        RECT 147.945 71.865 148.225 72.145 ;
        RECT 147.945 71.465 148.225 71.745 ;
        RECT 137.075 70.650 137.355 70.930 ;
        RECT 137.745 70.650 138.025 70.930 ;
        RECT 138.175 70.650 138.455 70.930 ;
        RECT 140.755 70.650 141.035 70.930 ;
        RECT 141.185 70.650 141.465 70.930 ;
        RECT 142.995 70.650 143.275 70.930 ;
        RECT 143.425 70.650 143.705 70.930 ;
        RECT 146.005 70.650 146.285 70.930 ;
        RECT 146.435 70.650 146.715 70.930 ;
        RECT 147.065 70.650 147.345 70.930 ;
        RECT 125.125 68.740 125.405 69.020 ;
        RECT 125.525 68.740 125.805 69.020 ;
        RECT 125.925 68.740 126.205 69.020 ;
        RECT 126.325 68.740 126.605 69.020 ;
        RECT 126.725 68.740 127.005 69.020 ;
        RECT 127.125 68.740 127.405 69.020 ;
        RECT 127.525 68.740 127.805 69.020 ;
        RECT 127.925 68.740 128.205 69.020 ;
        RECT 128.325 68.740 128.605 69.020 ;
        RECT 128.725 68.740 129.005 69.020 ;
        RECT 129.125 68.740 129.405 69.020 ;
        RECT 129.525 68.740 129.805 69.020 ;
        RECT 129.925 68.740 130.205 69.020 ;
        RECT 130.325 68.740 130.605 69.020 ;
        RECT 124.465 66.400 124.745 66.680 ;
        RECT 124.865 66.400 125.145 66.680 ;
        RECT 131.015 67.810 131.295 68.090 ;
        RECT 131.415 67.810 131.695 68.090 ;
        RECT 132.020 66.955 132.300 67.235 ;
        RECT 136.795 66.955 137.075 67.235 ;
        RECT 137.465 66.955 137.745 67.235 ;
        RECT 139.745 66.955 140.025 67.235 ;
        RECT 144.305 66.955 144.585 67.235 ;
        RECT 146.585 66.955 146.865 67.235 ;
        RECT 147.255 66.955 147.535 67.235 ;
        RECT 109.595 65.310 109.875 65.590 ;
        RECT 109.995 65.310 110.275 65.590 ;
        RECT 110.395 65.310 110.675 65.590 ;
        RECT 107.185 62.185 107.465 62.465 ;
        RECT 107.185 60.815 107.465 61.095 ;
        RECT 111.745 63.555 112.025 63.835 ;
        RECT 111.745 62.185 112.025 62.465 ;
        RECT 111.745 60.815 112.025 61.095 ;
        RECT 116.305 63.555 116.585 63.835 ;
        RECT 116.305 62.185 116.585 62.465 ;
        RECT 116.305 60.815 116.585 61.095 ;
        RECT 120.865 63.555 121.145 63.835 ;
        RECT 120.865 62.185 121.145 62.465 ;
        RECT 120.865 60.815 121.145 61.095 ;
        RECT 125.425 63.555 125.705 63.835 ;
        RECT 125.425 62.185 125.705 62.465 ;
        RECT 125.425 60.815 125.705 61.095 ;
        RECT 129.985 63.555 130.265 63.835 ;
        RECT 129.985 62.185 130.265 62.465 ;
        RECT 129.985 60.815 130.265 61.095 ;
        RECT 134.545 63.555 134.825 63.835 ;
        RECT 134.545 62.185 134.825 62.465 ;
        RECT 134.545 60.815 134.825 61.095 ;
        RECT 139.105 63.555 139.385 63.835 ;
        RECT 141.385 63.555 141.665 63.835 ;
        RECT 143.665 63.555 143.945 63.835 ;
        RECT 144.335 63.555 144.615 63.835 ;
        RECT 139.105 62.185 139.385 62.465 ;
        RECT 141.385 62.185 141.665 62.465 ;
        RECT 143.665 62.185 143.945 62.465 ;
        RECT 144.335 62.185 144.615 62.465 ;
        RECT 139.105 60.815 139.385 61.095 ;
        RECT 141.385 60.815 141.665 61.095 ;
        RECT 143.665 60.815 143.945 61.095 ;
        RECT 144.335 60.815 144.615 61.095 ;
        RECT 36.775 59.755 37.055 60.035 ;
        RECT 36.775 59.355 37.055 59.635 ;
        RECT 37.205 59.755 37.485 60.035 ;
        RECT 37.205 59.355 37.485 59.635 ;
        RECT 37.635 59.755 37.915 60.035 ;
        RECT 37.635 59.355 37.915 59.635 ;
        RECT 38.305 59.755 38.585 60.035 ;
        RECT 38.305 59.355 38.585 59.635 ;
        RECT 0.765 57.925 1.045 58.205 ;
        RECT 0.765 57.525 1.045 57.805 ;
        RECT 0.765 57.125 1.045 57.405 ;
        RECT 53.010 56.465 53.290 56.745 ;
        RECT 53.010 56.065 53.290 56.345 ;
        RECT 53.010 55.665 53.290 55.945 ;
        RECT 33.900 39.640 34.180 39.920 ;
        RECT 34.300 39.640 34.580 39.920 ;
        RECT 34.700 39.640 34.980 39.920 ;
        RECT 32.800 35.960 33.080 36.240 ;
        RECT 33.200 35.960 33.480 36.240 ;
        RECT 33.600 35.960 33.880 36.240 ;
        RECT 53.010 29.870 53.290 30.150 ;
        RECT 53.010 29.470 53.290 29.750 ;
        RECT 53.010 29.070 53.290 29.350 ;
        RECT 53.950 57.260 54.230 57.540 ;
        RECT 54.350 57.260 54.630 57.540 ;
        RECT 54.750 57.260 55.030 57.540 ;
        RECT 120.560 55.230 120.840 55.510 ;
        RECT 120.960 55.230 121.240 55.510 ;
        RECT 121.360 55.230 121.640 55.510 ;
        RECT 185.690 55.230 185.970 55.510 ;
        RECT 186.090 55.230 186.370 55.510 ;
        RECT 186.490 55.230 186.770 55.510 ;
        RECT 187.390 74.985 187.670 75.265 ;
        RECT 187.790 74.985 188.070 75.265 ;
        RECT 188.190 74.985 188.470 75.265 ;
        RECT 78.695 53.385 78.975 53.665 ;
        RECT 79.095 53.385 79.375 53.665 ;
        RECT 79.495 53.385 79.775 53.665 ;
        RECT 55.925 52.200 56.205 52.480 ;
        RECT 55.925 51.800 56.205 52.080 ;
        RECT 65.835 52.200 66.115 52.480 ;
        RECT 65.835 51.800 66.115 52.080 ;
        RECT 68.115 52.200 68.395 52.480 ;
        RECT 68.115 51.800 68.395 52.080 ;
        RECT 70.395 52.200 70.675 52.480 ;
        RECT 70.395 51.800 70.675 52.080 ;
        RECT 72.675 52.200 72.955 52.480 ;
        RECT 72.675 51.800 72.955 52.080 ;
        RECT 74.955 52.200 75.235 52.480 ;
        RECT 74.955 51.800 75.235 52.080 ;
        RECT 77.235 52.200 77.515 52.480 ;
        RECT 77.235 51.800 77.515 52.080 ;
        RECT 81.795 52.200 82.075 52.480 ;
        RECT 81.795 51.800 82.075 52.080 ;
        RECT 84.075 52.200 84.355 52.480 ;
        RECT 84.075 51.800 84.355 52.080 ;
        RECT 86.355 52.200 86.635 52.480 ;
        RECT 86.355 51.800 86.635 52.080 ;
        RECT 88.635 52.200 88.915 52.480 ;
        RECT 88.635 51.800 88.915 52.080 ;
        RECT 90.915 52.200 91.195 52.480 ;
        RECT 90.915 51.800 91.195 52.080 ;
        RECT 93.195 52.200 93.475 52.480 ;
        RECT 93.195 51.800 93.475 52.080 ;
        RECT 95.425 52.200 95.705 52.480 ;
        RECT 95.425 51.800 95.705 52.080 ;
        RECT 55.925 48.610 56.205 48.890 ;
        RECT 55.925 48.210 56.205 48.490 ;
        RECT 56.595 48.610 56.875 48.890 ;
        RECT 56.595 48.210 56.875 48.490 ;
        RECT 57.375 48.610 57.655 48.890 ;
        RECT 57.375 48.210 57.655 48.490 ;
        RECT 58.155 48.610 58.435 48.890 ;
        RECT 58.155 48.210 58.435 48.490 ;
        RECT 55.440 46.315 55.720 46.595 ;
        RECT 57.765 46.315 58.045 46.595 ;
        RECT 58.165 46.315 58.445 46.595 ;
        RECT 58.565 46.315 58.845 46.595 ;
        RECT 62.715 48.610 62.995 48.890 ;
        RECT 62.715 48.210 62.995 48.490 ;
        RECT 63.495 48.610 63.775 48.890 ;
        RECT 63.495 48.210 63.775 48.490 ;
        RECT 64.275 48.610 64.555 48.890 ;
        RECT 64.275 48.210 64.555 48.490 ;
        RECT 65.055 48.610 65.335 48.890 ;
        RECT 65.055 48.210 65.335 48.490 ;
        RECT 60.435 46.800 60.715 47.080 ;
        RECT 60.435 46.400 60.715 46.680 ;
        RECT 55.440 45.915 55.720 46.195 ;
        RECT 55.440 45.515 55.720 45.795 ;
        RECT 60.480 45.720 60.760 46.000 ;
        RECT 60.880 45.720 61.160 46.000 ;
        RECT 61.280 45.720 61.560 46.000 ;
        RECT 55.925 43.995 56.205 44.275 ;
        RECT 56.595 43.995 56.875 44.275 ;
        RECT 57.375 43.995 57.655 44.275 ;
        RECT 58.155 43.995 58.435 44.275 ;
        RECT 55.485 38.175 55.765 38.455 ;
        RECT 55.885 38.175 56.165 38.455 ;
        RECT 56.285 38.175 56.565 38.455 ;
        RECT 62.715 43.995 62.995 44.275 ;
        RECT 63.495 43.995 63.775 44.275 ;
        RECT 64.275 43.995 64.555 44.275 ;
        RECT 64.945 43.995 65.225 44.275 ;
        RECT 60.480 37.350 60.760 37.630 ;
        RECT 60.880 37.350 61.160 37.630 ;
        RECT 61.280 37.350 61.560 37.630 ;
        RECT 68.115 46.800 68.395 47.080 ;
        RECT 68.115 46.400 68.395 46.680 ;
        RECT 72.675 46.800 72.955 47.080 ;
        RECT 72.675 46.400 72.955 46.680 ;
        RECT 77.235 46.800 77.515 47.080 ;
        RECT 77.235 46.400 77.515 46.680 ;
        RECT 81.795 46.800 82.075 47.080 ;
        RECT 86.355 46.800 86.635 47.080 ;
        RECT 81.795 46.400 82.075 46.680 ;
        RECT 83.925 46.400 84.205 46.680 ;
        RECT 84.325 46.400 84.605 46.680 ;
        RECT 84.725 46.400 85.005 46.680 ;
        RECT 86.355 46.400 86.635 46.680 ;
        RECT 93.975 48.610 94.255 48.890 ;
        RECT 93.975 48.210 94.255 48.490 ;
        RECT 94.755 48.610 95.035 48.890 ;
        RECT 94.755 48.210 95.035 48.490 ;
        RECT 95.425 48.610 95.705 48.890 ;
        RECT 95.425 48.210 95.705 48.490 ;
        RECT 90.915 46.800 91.195 47.080 ;
        RECT 90.915 46.400 91.195 46.680 ;
        RECT 83.480 45.720 83.760 46.000 ;
        RECT 83.880 45.720 84.160 46.000 ;
        RECT 84.280 45.720 84.560 46.000 ;
        RECT 69.135 43.995 69.415 44.275 ;
        RECT 69.805 43.995 70.085 44.275 ;
        RECT 71.085 43.995 71.365 44.275 ;
        RECT 72.365 43.995 72.645 44.275 ;
        RECT 76.925 43.995 77.205 44.275 ;
        RECT 78.205 43.995 78.485 44.275 ;
        RECT 79.485 43.995 79.765 44.275 ;
        RECT 80.765 43.995 81.045 44.275 ;
        RECT 82.045 43.995 82.325 44.275 ;
        RECT 86.605 43.995 86.885 44.275 ;
        RECT 87.885 43.995 88.165 44.275 ;
        RECT 89.165 43.995 89.445 44.275 ;
        RECT 89.835 43.995 90.115 44.275 ;
        RECT 75.325 42.485 75.605 42.765 ;
        RECT 75.725 42.485 76.005 42.765 ;
        RECT 76.125 42.485 76.405 42.765 ;
        RECT 73.165 41.805 73.445 42.085 ;
        RECT 73.565 41.805 73.845 42.085 ;
        RECT 73.965 41.805 74.245 42.085 ;
        RECT 69.135 40.190 69.415 40.470 ;
        RECT 69.135 39.790 69.415 40.070 ;
        RECT 69.805 40.190 70.085 40.470 ;
        RECT 69.805 39.790 70.085 40.070 ;
        RECT 71.085 40.190 71.365 40.470 ;
        RECT 71.085 39.790 71.365 40.070 ;
        RECT 72.365 40.190 72.645 40.470 ;
        RECT 72.365 39.790 72.645 40.070 ;
        RECT 76.925 40.190 77.205 40.470 ;
        RECT 76.925 39.790 77.205 40.070 ;
        RECT 78.205 40.190 78.485 40.470 ;
        RECT 78.205 39.790 78.485 40.070 ;
        RECT 79.485 40.190 79.765 40.470 ;
        RECT 79.485 39.790 79.765 40.070 ;
        RECT 80.765 40.190 81.045 40.470 ;
        RECT 80.765 39.790 81.045 40.070 ;
        RECT 82.045 40.190 82.325 40.470 ;
        RECT 82.045 39.790 82.325 40.070 ;
        RECT 70.160 37.350 70.440 37.630 ;
        RECT 70.560 37.350 70.840 37.630 ;
        RECT 70.960 37.350 71.240 37.630 ;
        RECT 64.645 35.840 64.925 36.120 ;
        RECT 65.275 35.840 65.555 36.120 ;
        RECT 64.645 33.100 64.925 33.380 ;
        RECT 65.675 33.100 65.955 33.380 ;
        RECT 54.110 31.970 54.390 32.250 ;
        RECT 54.110 31.570 54.390 31.850 ;
        RECT 86.605 40.190 86.885 40.470 ;
        RECT 86.605 39.790 86.885 40.070 ;
        RECT 87.885 40.190 88.165 40.470 ;
        RECT 87.885 39.790 88.165 40.070 ;
        RECT 89.165 40.190 89.445 40.470 ;
        RECT 89.165 39.790 89.445 40.070 ;
        RECT 89.835 40.190 90.115 40.470 ;
        RECT 89.835 39.790 90.115 40.070 ;
        RECT 84.480 38.175 84.760 38.455 ;
        RECT 84.880 38.175 85.160 38.455 ;
        RECT 85.280 38.175 85.560 38.455 ;
        RECT 85.680 38.175 85.960 38.455 ;
        RECT 78.235 35.840 78.515 36.120 ;
        RECT 79.515 35.840 79.795 36.120 ;
        RECT 80.795 35.840 81.075 36.120 ;
        RECT 94.085 45.035 94.365 45.315 ;
        RECT 94.085 44.635 94.365 44.915 ;
        RECT 94.755 45.035 95.035 45.315 ;
        RECT 94.755 44.635 95.035 44.915 ;
        RECT 97.035 45.035 97.315 45.315 ;
        RECT 97.035 44.635 97.315 44.915 ;
        RECT 99.315 45.035 99.595 45.315 ;
        RECT 99.315 44.635 99.595 44.915 ;
        RECT 99.670 42.485 99.950 42.765 ;
        RECT 100.070 42.485 100.350 42.765 ;
        RECT 100.470 42.485 100.750 42.765 ;
        RECT 99.670 41.805 99.950 42.085 ;
        RECT 100.070 41.805 100.350 42.085 ;
        RECT 100.470 41.805 100.750 42.085 ;
        RECT 94.085 40.285 94.365 40.565 ;
        RECT 94.755 40.285 95.035 40.565 ;
        RECT 97.035 40.285 97.315 40.565 ;
        RECT 99.315 40.285 99.595 40.565 ;
        RECT 103.875 45.035 104.155 45.315 ;
        RECT 103.875 44.635 104.155 44.915 ;
        RECT 103.875 40.285 104.155 40.565 ;
        RECT 108.435 45.035 108.715 45.315 ;
        RECT 108.435 44.635 108.715 44.915 ;
        RECT 112.995 45.035 113.275 45.315 ;
        RECT 112.995 44.635 113.275 44.915 ;
        RECT 115.275 45.035 115.555 45.315 ;
        RECT 115.275 44.635 115.555 44.915 ;
        RECT 117.555 45.035 117.835 45.315 ;
        RECT 117.555 44.635 117.835 44.915 ;
        RECT 118.225 45.035 118.505 45.315 ;
        RECT 118.225 44.635 118.505 44.915 ;
        RECT 110.715 42.545 110.995 42.825 ;
        RECT 110.715 42.145 110.995 42.425 ;
        RECT 110.715 41.745 110.995 42.025 ;
        RECT 108.435 40.285 108.715 40.565 ;
        RECT 112.995 40.285 113.275 40.565 ;
        RECT 115.275 40.285 115.555 40.565 ;
        RECT 117.555 40.285 117.835 40.565 ;
        RECT 118.225 40.285 118.505 40.565 ;
        RECT 67.635 34.430 67.915 34.710 ;
        RECT 68.035 34.430 68.315 34.710 ;
        RECT 72.195 34.430 72.475 34.710 ;
        RECT 72.595 34.430 72.875 34.710 ;
        RECT 76.755 34.430 77.035 34.710 ;
        RECT 77.155 34.430 77.435 34.710 ;
        RECT 79.115 34.430 79.395 34.710 ;
        RECT 79.515 34.430 79.795 34.710 ;
        RECT 79.915 34.430 80.195 34.710 ;
        RECT 81.875 34.430 82.155 34.710 ;
        RECT 82.275 34.430 82.555 34.710 ;
        RECT 68.955 33.100 69.235 33.380 ;
        RECT 72.235 33.100 72.515 33.380 ;
        RECT 86.435 34.430 86.715 34.710 ;
        RECT 86.835 34.430 87.115 34.710 ;
        RECT 90.995 34.430 91.275 34.710 ;
        RECT 91.395 34.430 91.675 34.710 ;
        RECT 86.795 33.100 87.075 33.380 ;
        RECT 90.075 33.100 90.355 33.380 ;
        RECT 80.875 32.000 81.155 32.280 ;
        RECT 81.275 32.000 81.555 32.280 ;
        RECT 54.110 31.170 54.390 31.450 ;
        RECT 65.505 31.305 65.785 31.585 ;
        RECT 65.905 31.305 66.185 31.585 ;
        RECT 66.305 31.305 66.585 31.585 ;
        RECT 93.755 35.840 94.035 36.120 ;
        RECT 94.385 35.840 94.665 36.120 ;
        RECT 93.355 33.100 93.635 33.380 ;
        RECT 94.385 33.100 94.665 33.380 ;
        RECT 92.725 30.725 93.005 31.005 ;
        RECT 92.725 30.325 93.005 30.605 ;
        RECT 92.725 29.925 93.005 30.205 ;
        RECT 132.250 46.470 132.530 46.750 ;
        RECT 132.250 46.070 132.530 46.350 ;
        RECT 132.250 45.670 132.530 45.950 ;
        RECT 124.405 44.520 124.685 44.800 ;
        RECT 124.405 44.120 124.685 44.400 ;
        RECT 125.075 44.520 125.355 44.800 ;
        RECT 125.075 44.120 125.355 44.400 ;
        RECT 125.505 44.520 125.785 44.800 ;
        RECT 125.505 44.120 125.785 44.400 ;
        RECT 125.935 44.520 126.215 44.800 ;
        RECT 125.935 44.120 126.215 44.400 ;
        RECT 126.795 44.520 127.075 44.800 ;
        RECT 126.795 44.120 127.075 44.400 ;
        RECT 127.655 44.520 127.935 44.800 ;
        RECT 127.655 44.120 127.935 44.400 ;
        RECT 128.085 44.520 128.365 44.800 ;
        RECT 128.085 44.120 128.365 44.400 ;
        RECT 128.515 44.520 128.795 44.800 ;
        RECT 128.515 44.120 128.795 44.400 ;
        RECT 129.185 44.520 129.465 44.800 ;
        RECT 129.185 44.120 129.465 44.400 ;
        RECT 135.065 44.520 135.345 44.800 ;
        RECT 135.065 44.120 135.345 44.400 ;
        RECT 135.735 44.520 136.015 44.800 ;
        RECT 135.735 44.120 136.015 44.400 ;
        RECT 136.165 44.520 136.445 44.800 ;
        RECT 136.165 44.120 136.445 44.400 ;
        RECT 136.595 44.520 136.875 44.800 ;
        RECT 136.595 44.120 136.875 44.400 ;
        RECT 137.455 44.520 137.735 44.800 ;
        RECT 137.455 44.120 137.735 44.400 ;
        RECT 138.315 44.520 138.595 44.800 ;
        RECT 138.315 44.120 138.595 44.400 ;
        RECT 125.130 42.145 125.410 42.425 ;
        RECT 125.530 42.145 125.810 42.425 ;
        RECT 127.965 42.145 128.245 42.425 ;
        RECT 128.365 42.145 128.645 42.425 ;
        RECT 132.270 42.145 132.550 42.425 ;
        RECT 132.670 42.145 132.950 42.425 ;
        RECT 133.070 42.145 133.350 42.425 ;
        RECT 135.790 42.145 136.070 42.425 ;
        RECT 136.190 42.145 136.470 42.425 ;
        RECT 124.405 40.670 124.685 40.950 ;
        RECT 124.405 40.270 124.685 40.550 ;
        RECT 125.075 40.670 125.355 40.950 ;
        RECT 125.075 40.270 125.355 40.550 ;
        RECT 125.505 40.670 125.785 40.950 ;
        RECT 125.505 40.270 125.785 40.550 ;
        RECT 125.935 40.670 126.215 40.950 ;
        RECT 125.935 40.270 126.215 40.550 ;
        RECT 126.795 40.670 127.075 40.950 ;
        RECT 126.795 40.270 127.075 40.550 ;
        RECT 127.655 40.670 127.935 40.950 ;
        RECT 127.655 40.270 127.935 40.550 ;
        RECT 128.085 40.670 128.365 40.950 ;
        RECT 128.085 40.270 128.365 40.550 ;
        RECT 128.515 40.670 128.795 40.950 ;
        RECT 128.515 40.270 128.795 40.550 ;
        RECT 129.185 40.670 129.465 40.950 ;
        RECT 129.185 40.270 129.465 40.550 ;
        RECT 135.065 40.670 135.345 40.950 ;
        RECT 135.065 40.270 135.345 40.550 ;
        RECT 135.735 40.670 136.015 40.950 ;
        RECT 135.735 40.270 136.015 40.550 ;
        RECT 136.165 40.670 136.445 40.950 ;
        RECT 136.165 40.270 136.445 40.550 ;
        RECT 136.595 40.670 136.875 40.950 ;
        RECT 136.595 40.270 136.875 40.550 ;
        RECT 137.455 40.670 137.735 40.950 ;
        RECT 137.455 40.270 137.735 40.550 ;
        RECT 139.175 44.520 139.455 44.800 ;
        RECT 139.175 44.120 139.455 44.400 ;
        RECT 140.035 44.520 140.315 44.800 ;
        RECT 140.035 44.120 140.315 44.400 ;
        RECT 140.895 44.520 141.175 44.800 ;
        RECT 140.895 44.120 141.175 44.400 ;
        RECT 141.755 44.520 142.035 44.800 ;
        RECT 141.755 44.120 142.035 44.400 ;
        RECT 142.615 44.520 142.895 44.800 ;
        RECT 142.615 44.120 142.895 44.400 ;
        RECT 143.045 44.520 143.325 44.800 ;
        RECT 143.045 44.120 143.325 44.400 ;
        RECT 143.475 44.520 143.755 44.800 ;
        RECT 143.475 44.120 143.755 44.400 ;
        RECT 144.145 44.520 144.425 44.800 ;
        RECT 144.145 44.120 144.425 44.400 ;
        RECT 142.925 42.145 143.205 42.425 ;
        RECT 143.325 42.145 143.605 42.425 ;
        RECT 138.315 40.670 138.595 40.950 ;
        RECT 138.315 40.270 138.595 40.550 ;
        RECT 139.175 40.670 139.455 40.950 ;
        RECT 139.175 40.270 139.455 40.550 ;
        RECT 140.035 40.670 140.315 40.950 ;
        RECT 140.035 40.270 140.315 40.550 ;
        RECT 140.895 40.670 141.175 40.950 ;
        RECT 140.895 40.270 141.175 40.550 ;
        RECT 141.755 40.670 142.035 40.950 ;
        RECT 141.755 40.270 142.035 40.550 ;
        RECT 142.615 40.670 142.895 40.950 ;
        RECT 142.615 40.270 142.895 40.550 ;
        RECT 143.045 40.670 143.325 40.950 ;
        RECT 143.045 40.270 143.325 40.550 ;
        RECT 143.475 40.670 143.755 40.950 ;
        RECT 143.475 40.270 143.755 40.550 ;
        RECT 144.145 40.670 144.425 40.950 ;
        RECT 144.145 40.270 144.425 40.550 ;
        RECT 122.390 35.225 122.670 35.505 ;
        RECT 122.390 34.825 122.670 35.105 ;
        RECT 123.520 38.110 123.800 38.390 ;
        RECT 129.170 38.110 129.450 38.390 ;
        RECT 129.570 38.110 129.850 38.390 ;
        RECT 129.970 38.110 130.250 38.390 ;
        RECT 123.520 37.710 123.800 37.990 ;
        RECT 123.520 37.310 123.800 37.590 ;
        RECT 120.720 30.990 121.000 31.270 ;
        RECT 120.720 30.590 121.000 30.870 ;
        RECT 120.720 30.190 121.000 30.470 ;
        RECT 65.505 29.205 65.785 29.485 ;
        RECT 65.905 29.205 66.185 29.485 ;
        RECT 66.305 29.205 66.585 29.485 ;
        RECT 64.645 27.410 64.925 27.690 ;
        RECT 65.675 27.410 65.955 27.690 ;
        RECT 64.645 24.670 64.925 24.950 ;
        RECT 65.275 24.670 65.555 24.950 ;
        RECT 80.875 28.510 81.155 28.790 ;
        RECT 81.275 28.510 81.555 28.790 ;
        RECT 68.955 27.410 69.235 27.690 ;
        RECT 72.235 27.410 72.515 27.690 ;
        RECT 67.635 26.080 67.915 26.360 ;
        RECT 68.035 26.080 68.315 26.360 ;
        RECT 72.195 26.080 72.475 26.360 ;
        RECT 72.595 26.080 72.875 26.360 ;
        RECT 86.795 27.410 87.075 27.690 ;
        RECT 90.075 27.410 90.355 27.690 ;
        RECT 76.755 26.080 77.035 26.360 ;
        RECT 77.155 26.080 77.435 26.360 ;
        RECT 79.115 26.080 79.395 26.360 ;
        RECT 79.515 26.080 79.795 26.360 ;
        RECT 79.915 26.080 80.195 26.360 ;
        RECT 81.875 26.080 82.155 26.360 ;
        RECT 82.275 26.080 82.555 26.360 ;
        RECT 86.435 26.080 86.715 26.360 ;
        RECT 86.835 26.080 87.115 26.360 ;
        RECT 90.995 26.080 91.275 26.360 ;
        RECT 91.395 26.080 91.675 26.360 ;
        RECT 60.480 23.160 60.760 23.440 ;
        RECT 60.880 23.160 61.160 23.440 ;
        RECT 61.280 23.160 61.560 23.440 ;
        RECT 55.485 22.335 55.765 22.615 ;
        RECT 55.885 22.335 56.165 22.615 ;
        RECT 56.285 22.335 56.565 22.615 ;
        RECT 55.925 16.515 56.205 16.795 ;
        RECT 56.595 16.515 56.875 16.795 ;
        RECT 57.375 16.515 57.655 16.795 ;
        RECT 58.155 16.515 58.435 16.795 ;
        RECT 62.715 16.515 62.995 16.795 ;
        RECT 63.495 16.515 63.775 16.795 ;
        RECT 64.275 16.515 64.555 16.795 ;
        RECT 64.945 16.515 65.225 16.795 ;
        RECT 55.440 14.995 55.720 15.275 ;
        RECT 55.440 14.595 55.720 14.875 ;
        RECT 60.480 14.790 60.760 15.070 ;
        RECT 60.880 14.790 61.160 15.070 ;
        RECT 61.280 14.790 61.560 15.070 ;
        RECT 55.440 14.195 55.720 14.475 ;
        RECT 57.765 14.195 58.045 14.475 ;
        RECT 58.165 14.195 58.445 14.475 ;
        RECT 58.565 14.195 58.845 14.475 ;
        RECT 60.435 14.110 60.715 14.390 ;
        RECT 60.435 13.710 60.715 13.990 ;
        RECT 55.925 12.300 56.205 12.580 ;
        RECT 55.925 11.900 56.205 12.180 ;
        RECT 56.595 12.300 56.875 12.580 ;
        RECT 56.595 11.900 56.875 12.180 ;
        RECT 57.375 12.300 57.655 12.580 ;
        RECT 57.375 11.900 57.655 12.180 ;
        RECT 58.155 12.300 58.435 12.580 ;
        RECT 58.155 11.900 58.435 12.180 ;
        RECT 78.235 24.670 78.515 24.950 ;
        RECT 79.515 24.670 79.795 24.950 ;
        RECT 80.795 24.670 81.075 24.950 ;
        RECT 70.160 23.160 70.440 23.440 ;
        RECT 70.560 23.160 70.840 23.440 ;
        RECT 70.960 23.160 71.240 23.440 ;
        RECT 69.135 20.720 69.415 21.000 ;
        RECT 69.135 20.320 69.415 20.600 ;
        RECT 69.805 20.720 70.085 21.000 ;
        RECT 69.805 20.320 70.085 20.600 ;
        RECT 71.085 20.720 71.365 21.000 ;
        RECT 71.085 20.320 71.365 20.600 ;
        RECT 72.365 20.720 72.645 21.000 ;
        RECT 72.365 20.320 72.645 20.600 ;
        RECT 93.355 27.410 93.635 27.690 ;
        RECT 94.385 27.410 94.665 27.690 ;
        RECT 124.170 37.330 124.450 37.610 ;
        RECT 124.570 37.330 124.850 37.610 ;
        RECT 124.970 37.330 125.250 37.610 ;
        RECT 126.515 37.330 126.795 37.610 ;
        RECT 126.915 37.330 127.195 37.610 ;
        RECT 124.755 36.600 125.035 36.880 ;
        RECT 124.755 36.200 125.035 36.480 ;
        RECT 125.425 36.600 125.705 36.880 ;
        RECT 125.425 36.200 125.705 36.480 ;
        RECT 125.855 36.600 126.135 36.880 ;
        RECT 125.855 36.200 126.135 36.480 ;
        RECT 126.285 36.600 126.565 36.880 ;
        RECT 126.285 36.200 126.565 36.480 ;
        RECT 127.145 36.600 127.425 36.880 ;
        RECT 127.145 36.200 127.425 36.480 ;
        RECT 128.005 36.600 128.285 36.880 ;
        RECT 128.005 36.200 128.285 36.480 ;
        RECT 128.435 36.600 128.715 36.880 ;
        RECT 128.435 36.200 128.715 36.480 ;
        RECT 128.865 36.600 129.145 36.880 ;
        RECT 128.865 36.200 129.145 36.480 ;
        RECT 129.515 36.600 129.795 36.880 ;
        RECT 129.515 36.200 129.795 36.480 ;
        RECT 135.065 36.700 135.345 36.980 ;
        RECT 135.065 36.300 135.345 36.580 ;
        RECT 135.735 36.700 136.015 36.980 ;
        RECT 135.735 36.300 136.015 36.580 ;
        RECT 136.165 36.700 136.445 36.980 ;
        RECT 136.165 36.300 136.445 36.580 ;
        RECT 136.595 36.700 136.875 36.980 ;
        RECT 136.595 36.300 136.875 36.580 ;
        RECT 137.455 36.700 137.735 36.980 ;
        RECT 137.455 36.300 137.735 36.580 ;
        RECT 138.315 36.700 138.595 36.980 ;
        RECT 138.315 36.300 138.595 36.580 ;
        RECT 125.595 34.825 125.875 35.105 ;
        RECT 125.995 34.825 126.275 35.105 ;
        RECT 128.215 34.825 128.495 35.105 ;
        RECT 128.615 34.825 128.895 35.105 ;
        RECT 129.170 34.825 129.450 35.105 ;
        RECT 129.570 34.825 129.850 35.105 ;
        RECT 129.970 34.825 130.250 35.105 ;
        RECT 135.790 34.825 136.070 35.105 ;
        RECT 136.190 34.825 136.470 35.105 ;
        RECT 124.755 33.375 125.035 33.655 ;
        RECT 124.755 32.975 125.035 33.255 ;
        RECT 125.425 33.375 125.705 33.655 ;
        RECT 125.425 32.975 125.705 33.255 ;
        RECT 125.855 33.375 126.135 33.655 ;
        RECT 125.855 32.975 126.135 33.255 ;
        RECT 128.435 33.375 128.715 33.655 ;
        RECT 128.435 32.975 128.715 33.255 ;
        RECT 128.865 33.375 129.145 33.655 ;
        RECT 128.865 32.975 129.145 33.255 ;
        RECT 129.515 33.375 129.795 33.655 ;
        RECT 129.515 32.975 129.795 33.255 ;
        RECT 135.065 32.850 135.345 33.130 ;
        RECT 135.065 32.450 135.345 32.730 ;
        RECT 124.755 31.800 125.035 32.080 ;
        RECT 124.755 31.400 125.035 31.680 ;
        RECT 125.425 31.800 125.705 32.080 ;
        RECT 125.425 31.400 125.705 31.680 ;
        RECT 125.855 31.800 126.135 32.080 ;
        RECT 125.855 31.400 126.135 31.680 ;
        RECT 126.285 31.800 126.565 32.080 ;
        RECT 126.285 31.400 126.565 31.680 ;
        RECT 127.145 31.800 127.425 32.080 ;
        RECT 127.145 31.400 127.425 31.680 ;
        RECT 135.735 32.850 136.015 33.130 ;
        RECT 135.735 32.450 136.015 32.730 ;
        RECT 136.165 32.850 136.445 33.130 ;
        RECT 136.165 32.450 136.445 32.730 ;
        RECT 136.595 32.850 136.875 33.130 ;
        RECT 136.595 32.450 136.875 32.730 ;
        RECT 128.005 31.800 128.285 32.080 ;
        RECT 128.005 31.400 128.285 31.680 ;
        RECT 128.435 31.800 128.715 32.080 ;
        RECT 128.435 31.400 128.715 31.680 ;
        RECT 128.865 31.800 129.145 32.080 ;
        RECT 128.865 31.400 129.145 31.680 ;
        RECT 129.515 31.800 129.795 32.080 ;
        RECT 137.455 32.850 137.735 33.130 ;
        RECT 137.455 32.450 137.735 32.730 ;
        RECT 139.175 36.700 139.455 36.980 ;
        RECT 139.175 36.300 139.455 36.580 ;
        RECT 140.035 36.700 140.315 36.980 ;
        RECT 140.035 36.300 140.315 36.580 ;
        RECT 140.895 36.700 141.175 36.980 ;
        RECT 140.895 36.300 141.175 36.580 ;
        RECT 141.755 36.700 142.035 36.980 ;
        RECT 141.755 36.300 142.035 36.580 ;
        RECT 142.615 36.700 142.895 36.980 ;
        RECT 142.615 36.300 142.895 36.580 ;
        RECT 143.045 36.700 143.325 36.980 ;
        RECT 143.045 36.300 143.325 36.580 ;
        RECT 143.475 36.700 143.755 36.980 ;
        RECT 143.475 36.300 143.755 36.580 ;
        RECT 144.145 36.700 144.425 36.980 ;
        RECT 144.145 36.300 144.425 36.580 ;
        RECT 142.925 34.825 143.205 35.105 ;
        RECT 143.325 34.825 143.605 35.105 ;
        RECT 138.315 32.850 138.595 33.130 ;
        RECT 138.315 32.450 138.595 32.730 ;
        RECT 139.175 32.850 139.455 33.130 ;
        RECT 139.175 32.450 139.455 32.730 ;
        RECT 140.035 32.850 140.315 33.130 ;
        RECT 140.035 32.450 140.315 32.730 ;
        RECT 140.895 32.850 141.175 33.130 ;
        RECT 140.895 32.450 141.175 32.730 ;
        RECT 141.755 32.850 142.035 33.130 ;
        RECT 141.755 32.450 142.035 32.730 ;
        RECT 142.615 32.850 142.895 33.130 ;
        RECT 142.615 32.450 142.895 32.730 ;
        RECT 143.045 32.850 143.325 33.130 ;
        RECT 143.045 32.450 143.325 32.730 ;
        RECT 143.475 32.850 143.755 33.130 ;
        RECT 143.475 32.450 143.755 32.730 ;
        RECT 144.145 32.850 144.425 33.130 ;
        RECT 144.145 32.450 144.425 32.730 ;
        RECT 129.515 31.400 129.795 31.680 ;
        RECT 124.170 30.670 124.450 30.950 ;
        RECT 124.570 30.670 124.850 30.950 ;
        RECT 124.970 30.670 125.250 30.950 ;
        RECT 126.745 30.670 127.025 30.950 ;
        RECT 127.145 30.670 127.425 30.950 ;
        RECT 127.545 30.670 127.825 30.950 ;
        RECT 129.990 30.670 130.270 30.950 ;
        RECT 129.990 30.270 130.270 30.550 ;
        RECT 123.520 26.255 123.800 26.535 ;
        RECT 123.520 25.855 123.800 26.135 ;
        RECT 123.520 25.455 123.800 25.735 ;
        RECT 124.170 29.610 124.450 29.890 ;
        RECT 124.570 29.610 124.850 29.890 ;
        RECT 124.970 29.610 125.250 29.890 ;
        RECT 126.745 29.610 127.025 29.890 ;
        RECT 127.145 29.610 127.425 29.890 ;
        RECT 127.545 29.610 127.825 29.890 ;
        RECT 129.990 29.870 130.270 30.150 ;
        RECT 93.755 24.670 94.035 24.950 ;
        RECT 94.385 24.670 94.665 24.950 ;
        RECT 84.480 22.335 84.760 22.615 ;
        RECT 84.880 22.335 85.160 22.615 ;
        RECT 85.280 22.335 85.560 22.615 ;
        RECT 85.680 22.335 85.960 22.615 ;
        RECT 76.925 20.720 77.205 21.000 ;
        RECT 76.925 20.320 77.205 20.600 ;
        RECT 78.205 20.720 78.485 21.000 ;
        RECT 78.205 20.320 78.485 20.600 ;
        RECT 79.485 20.720 79.765 21.000 ;
        RECT 79.485 20.320 79.765 20.600 ;
        RECT 80.765 20.720 81.045 21.000 ;
        RECT 80.765 20.320 81.045 20.600 ;
        RECT 82.045 20.720 82.325 21.000 ;
        RECT 82.045 20.320 82.325 20.600 ;
        RECT 86.605 20.720 86.885 21.000 ;
        RECT 86.605 20.320 86.885 20.600 ;
        RECT 87.885 20.720 88.165 21.000 ;
        RECT 87.885 20.320 88.165 20.600 ;
        RECT 89.165 20.720 89.445 21.000 ;
        RECT 89.165 20.320 89.445 20.600 ;
        RECT 89.835 20.720 90.115 21.000 ;
        RECT 89.835 20.320 90.115 20.600 ;
        RECT 73.165 18.705 73.445 18.985 ;
        RECT 73.565 18.705 73.845 18.985 ;
        RECT 73.965 18.705 74.245 18.985 ;
        RECT 75.325 18.025 75.605 18.305 ;
        RECT 75.725 18.025 76.005 18.305 ;
        RECT 76.125 18.025 76.405 18.305 ;
        RECT 69.135 16.515 69.415 16.795 ;
        RECT 69.805 16.515 70.085 16.795 ;
        RECT 71.085 16.515 71.365 16.795 ;
        RECT 72.365 16.515 72.645 16.795 ;
        RECT 76.925 16.515 77.205 16.795 ;
        RECT 78.205 16.515 78.485 16.795 ;
        RECT 79.485 16.515 79.765 16.795 ;
        RECT 80.765 16.515 81.045 16.795 ;
        RECT 82.045 16.515 82.325 16.795 ;
        RECT 86.605 16.515 86.885 16.795 ;
        RECT 87.885 16.515 88.165 16.795 ;
        RECT 89.165 16.515 89.445 16.795 ;
        RECT 89.835 16.515 90.115 16.795 ;
        RECT 68.115 14.110 68.395 14.390 ;
        RECT 68.115 13.710 68.395 13.990 ;
        RECT 62.715 12.300 62.995 12.580 ;
        RECT 62.715 11.900 62.995 12.180 ;
        RECT 63.495 12.300 63.775 12.580 ;
        RECT 63.495 11.900 63.775 12.180 ;
        RECT 64.275 12.300 64.555 12.580 ;
        RECT 64.275 11.900 64.555 12.180 ;
        RECT 65.055 12.300 65.335 12.580 ;
        RECT 65.055 11.900 65.335 12.180 ;
        RECT 83.480 14.790 83.760 15.070 ;
        RECT 83.880 14.790 84.160 15.070 ;
        RECT 84.280 14.790 84.560 15.070 ;
        RECT 72.675 14.110 72.955 14.390 ;
        RECT 72.675 13.710 72.955 13.990 ;
        RECT 77.235 14.110 77.515 14.390 ;
        RECT 77.235 13.710 77.515 13.990 ;
        RECT 81.795 14.110 82.075 14.390 ;
        RECT 83.925 14.110 84.205 14.390 ;
        RECT 84.325 14.110 84.605 14.390 ;
        RECT 84.725 14.110 85.005 14.390 ;
        RECT 86.355 14.110 86.635 14.390 ;
        RECT 81.795 13.710 82.075 13.990 ;
        RECT 86.355 13.710 86.635 13.990 ;
        RECT 90.915 14.110 91.195 14.390 ;
        RECT 90.915 13.710 91.195 13.990 ;
        RECT 124.755 28.880 125.035 29.160 ;
        RECT 124.755 28.480 125.035 28.760 ;
        RECT 125.425 28.880 125.705 29.160 ;
        RECT 125.425 28.480 125.705 28.760 ;
        RECT 125.855 28.880 126.135 29.160 ;
        RECT 125.855 28.480 126.135 28.760 ;
        RECT 126.285 28.880 126.565 29.160 ;
        RECT 126.285 28.480 126.565 28.760 ;
        RECT 127.145 28.880 127.425 29.160 ;
        RECT 127.145 28.480 127.425 28.760 ;
        RECT 128.005 28.880 128.285 29.160 ;
        RECT 128.005 28.480 128.285 28.760 ;
        RECT 128.435 28.880 128.715 29.160 ;
        RECT 128.435 28.480 128.715 28.760 ;
        RECT 128.865 28.880 129.145 29.160 ;
        RECT 128.865 28.480 129.145 28.760 ;
        RECT 129.515 28.880 129.795 29.160 ;
        RECT 129.515 28.480 129.795 28.760 ;
        RECT 124.755 27.305 125.035 27.585 ;
        RECT 124.755 26.905 125.035 27.185 ;
        RECT 125.425 27.305 125.705 27.585 ;
        RECT 125.425 26.905 125.705 27.185 ;
        RECT 125.855 27.305 126.135 27.585 ;
        RECT 125.855 26.905 126.135 27.185 ;
        RECT 135.065 29.760 135.345 30.040 ;
        RECT 135.065 29.360 135.345 29.640 ;
        RECT 135.735 29.760 136.015 30.040 ;
        RECT 135.735 29.360 136.015 29.640 ;
        RECT 136.165 29.760 136.445 30.040 ;
        RECT 136.165 29.360 136.445 29.640 ;
        RECT 136.595 29.760 136.875 30.040 ;
        RECT 136.595 29.360 136.875 29.640 ;
        RECT 137.455 29.760 137.735 30.040 ;
        RECT 137.455 29.360 137.735 29.640 ;
        RECT 138.315 29.760 138.595 30.040 ;
        RECT 138.315 29.360 138.595 29.640 ;
        RECT 128.435 27.305 128.715 27.585 ;
        RECT 128.435 26.905 128.715 27.185 ;
        RECT 128.865 27.305 129.145 27.585 ;
        RECT 128.865 26.905 129.145 27.185 ;
        RECT 129.515 27.305 129.795 27.585 ;
        RECT 129.515 26.905 129.795 27.185 ;
        RECT 131.200 27.385 131.480 27.665 ;
        RECT 131.600 27.385 131.880 27.665 ;
        RECT 135.790 27.385 136.070 27.665 ;
        RECT 136.190 27.385 136.470 27.665 ;
        RECT 125.595 25.455 125.875 25.735 ;
        RECT 125.995 25.455 126.275 25.735 ;
        RECT 128.215 25.455 128.495 25.735 ;
        RECT 128.615 25.455 128.895 25.735 ;
        RECT 129.170 25.455 129.450 25.735 ;
        RECT 129.570 25.455 129.850 25.735 ;
        RECT 129.970 25.455 130.250 25.735 ;
        RECT 135.065 25.910 135.345 26.190 ;
        RECT 135.065 25.510 135.345 25.790 ;
        RECT 124.755 24.080 125.035 24.360 ;
        RECT 124.755 23.680 125.035 23.960 ;
        RECT 125.425 24.080 125.705 24.360 ;
        RECT 125.425 23.680 125.705 23.960 ;
        RECT 125.855 24.080 126.135 24.360 ;
        RECT 125.855 23.680 126.135 23.960 ;
        RECT 126.285 24.080 126.565 24.360 ;
        RECT 126.285 23.680 126.565 23.960 ;
        RECT 127.145 24.080 127.425 24.360 ;
        RECT 127.145 23.680 127.425 23.960 ;
        RECT 135.735 25.910 136.015 26.190 ;
        RECT 135.735 25.510 136.015 25.790 ;
        RECT 136.165 25.910 136.445 26.190 ;
        RECT 136.165 25.510 136.445 25.790 ;
        RECT 136.595 25.910 136.875 26.190 ;
        RECT 136.595 25.510 136.875 25.790 ;
        RECT 137.455 25.910 137.735 26.190 ;
        RECT 137.455 25.510 137.735 25.790 ;
        RECT 139.175 29.760 139.455 30.040 ;
        RECT 139.175 29.360 139.455 29.640 ;
        RECT 140.035 29.760 140.315 30.040 ;
        RECT 140.035 29.360 140.315 29.640 ;
        RECT 140.895 29.760 141.175 30.040 ;
        RECT 140.895 29.360 141.175 29.640 ;
        RECT 141.755 29.760 142.035 30.040 ;
        RECT 141.755 29.360 142.035 29.640 ;
        RECT 142.615 29.760 142.895 30.040 ;
        RECT 142.615 29.360 142.895 29.640 ;
        RECT 143.045 29.760 143.325 30.040 ;
        RECT 143.045 29.360 143.325 29.640 ;
        RECT 143.475 29.760 143.755 30.040 ;
        RECT 143.475 29.360 143.755 29.640 ;
        RECT 144.145 29.760 144.425 30.040 ;
        RECT 144.145 29.360 144.425 29.640 ;
        RECT 142.925 27.385 143.205 27.665 ;
        RECT 143.325 27.385 143.605 27.665 ;
        RECT 138.315 25.910 138.595 26.190 ;
        RECT 138.315 25.510 138.595 25.790 ;
        RECT 139.175 25.910 139.455 26.190 ;
        RECT 139.175 25.510 139.455 25.790 ;
        RECT 140.035 25.910 140.315 26.190 ;
        RECT 140.035 25.510 140.315 25.790 ;
        RECT 140.895 25.910 141.175 26.190 ;
        RECT 140.895 25.510 141.175 25.790 ;
        RECT 141.755 25.910 142.035 26.190 ;
        RECT 141.755 25.510 142.035 25.790 ;
        RECT 142.615 25.910 142.895 26.190 ;
        RECT 142.615 25.510 142.895 25.790 ;
        RECT 143.045 25.910 143.325 26.190 ;
        RECT 143.045 25.510 143.325 25.790 ;
        RECT 143.475 25.910 143.755 26.190 ;
        RECT 143.475 25.510 143.755 25.790 ;
        RECT 144.145 25.910 144.425 26.190 ;
        RECT 144.145 25.510 144.425 25.790 ;
        RECT 128.005 24.080 128.285 24.360 ;
        RECT 128.005 23.680 128.285 23.960 ;
        RECT 128.435 24.080 128.715 24.360 ;
        RECT 128.435 23.680 128.715 23.960 ;
        RECT 128.865 24.080 129.145 24.360 ;
        RECT 128.865 23.680 129.145 23.960 ;
        RECT 129.515 24.080 129.795 24.360 ;
        RECT 129.515 23.680 129.795 23.960 ;
        RECT 188.200 74.050 188.480 74.330 ;
        RECT 188.200 73.650 188.480 73.930 ;
        RECT 188.200 73.250 188.480 73.530 ;
        RECT 203.130 86.705 203.410 86.985 ;
        RECT 203.130 86.305 203.410 86.585 ;
        RECT 203.130 85.905 203.410 86.185 ;
        RECT 203.130 85.505 203.410 85.785 ;
        RECT 194.365 69.540 194.645 69.820 ;
        RECT 194.365 69.140 194.645 69.420 ;
        RECT 189.165 68.740 189.445 69.020 ;
        RECT 194.365 68.740 194.645 69.020 ;
        RECT 189.165 68.340 189.445 68.620 ;
        RECT 189.165 67.940 189.445 68.220 ;
        RECT 189.165 56.995 189.445 57.275 ;
        RECT 189.165 56.595 189.445 56.875 ;
        RECT 189.165 56.195 189.445 56.475 ;
        RECT 199.710 63.495 199.990 63.775 ;
        RECT 199.710 63.095 199.990 63.375 ;
        RECT 190.690 42.145 190.970 42.425 ;
        RECT 191.090 42.145 191.370 42.425 ;
        RECT 191.490 42.145 191.770 42.425 ;
        RECT 188.200 39.360 188.480 39.640 ;
        RECT 188.200 38.960 188.480 39.240 ;
        RECT 188.200 38.560 188.480 38.840 ;
        RECT 186.550 23.305 186.830 23.585 ;
        RECT 186.950 23.305 187.230 23.585 ;
        RECT 187.350 23.305 187.630 23.585 ;
        RECT 124.170 22.950 124.450 23.230 ;
        RECT 124.570 22.950 124.850 23.230 ;
        RECT 124.970 22.950 125.250 23.230 ;
        RECT 126.515 22.950 126.795 23.230 ;
        RECT 126.915 22.950 127.195 23.230 ;
        RECT 135.065 20.740 135.345 21.020 ;
        RECT 94.085 20.225 94.365 20.505 ;
        RECT 94.755 20.225 95.035 20.505 ;
        RECT 97.035 20.225 97.315 20.505 ;
        RECT 99.315 20.225 99.595 20.505 ;
        RECT 99.670 18.705 99.950 18.985 ;
        RECT 100.070 18.705 100.350 18.985 ;
        RECT 100.470 18.705 100.750 18.985 ;
        RECT 99.670 18.025 99.950 18.305 ;
        RECT 100.070 18.025 100.350 18.305 ;
        RECT 100.470 18.025 100.750 18.305 ;
        RECT 94.085 15.875 94.365 16.155 ;
        RECT 94.085 15.475 94.365 15.755 ;
        RECT 94.755 15.875 95.035 16.155 ;
        RECT 94.755 15.475 95.035 15.755 ;
        RECT 97.035 15.875 97.315 16.155 ;
        RECT 97.035 15.475 97.315 15.755 ;
        RECT 99.315 15.875 99.595 16.155 ;
        RECT 99.315 15.475 99.595 15.755 ;
        RECT 103.875 20.225 104.155 20.505 ;
        RECT 103.875 15.875 104.155 16.155 ;
        RECT 103.875 15.475 104.155 15.755 ;
        RECT 108.435 20.225 108.715 20.505 ;
        RECT 112.995 20.225 113.275 20.505 ;
        RECT 115.275 20.225 115.555 20.505 ;
        RECT 117.555 20.225 117.835 20.505 ;
        RECT 118.225 20.225 118.505 20.505 ;
        RECT 135.065 20.340 135.345 20.620 ;
        RECT 135.735 20.740 136.015 21.020 ;
        RECT 135.735 20.340 136.015 20.620 ;
        RECT 136.165 20.740 136.445 21.020 ;
        RECT 136.165 20.340 136.445 20.620 ;
        RECT 136.595 20.740 136.875 21.020 ;
        RECT 136.595 20.340 136.875 20.620 ;
        RECT 110.715 18.765 110.995 19.045 ;
        RECT 137.455 20.740 137.735 21.020 ;
        RECT 137.455 20.340 137.735 20.620 ;
        RECT 138.315 20.740 138.595 21.020 ;
        RECT 138.315 20.340 138.595 20.620 ;
        RECT 110.715 18.365 110.995 18.645 ;
        RECT 135.790 18.365 136.070 18.645 ;
        RECT 136.190 18.365 136.470 18.645 ;
        RECT 110.715 17.965 110.995 18.245 ;
        RECT 108.435 15.875 108.715 16.155 ;
        RECT 108.435 15.475 108.715 15.755 ;
        RECT 135.065 16.890 135.345 17.170 ;
        RECT 135.065 16.490 135.345 16.770 ;
        RECT 135.735 16.890 136.015 17.170 ;
        RECT 135.735 16.490 136.015 16.770 ;
        RECT 136.165 16.890 136.445 17.170 ;
        RECT 136.165 16.490 136.445 16.770 ;
        RECT 136.595 16.890 136.875 17.170 ;
        RECT 136.595 16.490 136.875 16.770 ;
        RECT 137.455 16.890 137.735 17.170 ;
        RECT 137.455 16.490 137.735 16.770 ;
        RECT 139.175 20.740 139.455 21.020 ;
        RECT 139.175 20.340 139.455 20.620 ;
        RECT 140.035 20.740 140.315 21.020 ;
        RECT 140.035 20.340 140.315 20.620 ;
        RECT 140.895 20.740 141.175 21.020 ;
        RECT 140.895 20.340 141.175 20.620 ;
        RECT 141.755 20.740 142.035 21.020 ;
        RECT 141.755 20.340 142.035 20.620 ;
        RECT 142.615 20.740 142.895 21.020 ;
        RECT 142.615 20.340 142.895 20.620 ;
        RECT 143.045 20.740 143.325 21.020 ;
        RECT 143.045 20.340 143.325 20.620 ;
        RECT 143.475 20.740 143.755 21.020 ;
        RECT 143.475 20.340 143.755 20.620 ;
        RECT 144.145 20.740 144.425 21.020 ;
        RECT 144.145 20.340 144.425 20.620 ;
        RECT 142.925 18.365 143.205 18.645 ;
        RECT 143.325 18.365 143.605 18.645 ;
        RECT 138.315 16.890 138.595 17.170 ;
        RECT 138.315 16.490 138.595 16.770 ;
        RECT 139.175 16.890 139.455 17.170 ;
        RECT 139.175 16.490 139.455 16.770 ;
        RECT 140.035 16.890 140.315 17.170 ;
        RECT 140.035 16.490 140.315 16.770 ;
        RECT 140.895 16.890 141.175 17.170 ;
        RECT 140.895 16.490 141.175 16.770 ;
        RECT 141.755 16.890 142.035 17.170 ;
        RECT 141.755 16.490 142.035 16.770 ;
        RECT 142.615 16.890 142.895 17.170 ;
        RECT 142.615 16.490 142.895 16.770 ;
        RECT 143.045 16.890 143.325 17.170 ;
        RECT 143.045 16.490 143.325 16.770 ;
        RECT 143.475 16.890 143.755 17.170 ;
        RECT 143.475 16.490 143.755 16.770 ;
        RECT 144.145 16.890 144.425 17.170 ;
        RECT 144.145 16.490 144.425 16.770 ;
        RECT 112.995 15.875 113.275 16.155 ;
        RECT 112.995 15.475 113.275 15.755 ;
        RECT 115.275 15.875 115.555 16.155 ;
        RECT 115.275 15.475 115.555 15.755 ;
        RECT 117.555 15.875 117.835 16.155 ;
        RECT 117.555 15.475 117.835 15.755 ;
        RECT 118.225 15.875 118.505 16.155 ;
        RECT 118.225 15.475 118.505 15.755 ;
        RECT 93.975 12.300 94.255 12.580 ;
        RECT 93.975 11.900 94.255 12.180 ;
        RECT 94.755 12.300 95.035 12.580 ;
        RECT 94.755 11.900 95.035 12.180 ;
        RECT 95.425 12.300 95.705 12.580 ;
        RECT 95.425 11.900 95.705 12.180 ;
        RECT 55.925 8.710 56.205 8.990 ;
        RECT 55.925 8.310 56.205 8.590 ;
        RECT 65.835 8.710 66.115 8.990 ;
        RECT 65.835 8.310 66.115 8.590 ;
        RECT 68.115 8.710 68.395 8.990 ;
        RECT 68.115 8.310 68.395 8.590 ;
        RECT 70.395 8.710 70.675 8.990 ;
        RECT 70.395 8.310 70.675 8.590 ;
        RECT 72.675 8.710 72.955 8.990 ;
        RECT 72.675 8.310 72.955 8.590 ;
        RECT 74.955 8.710 75.235 8.990 ;
        RECT 74.955 8.310 75.235 8.590 ;
        RECT 77.235 8.710 77.515 8.990 ;
        RECT 77.235 8.310 77.515 8.590 ;
        RECT 81.795 8.710 82.075 8.990 ;
        RECT 81.795 8.310 82.075 8.590 ;
        RECT 84.075 8.710 84.355 8.990 ;
        RECT 84.075 8.310 84.355 8.590 ;
        RECT 86.355 8.710 86.635 8.990 ;
        RECT 86.355 8.310 86.635 8.590 ;
        RECT 88.635 8.710 88.915 8.990 ;
        RECT 88.635 8.310 88.915 8.590 ;
        RECT 90.915 8.710 91.195 8.990 ;
        RECT 90.915 8.310 91.195 8.590 ;
        RECT 93.195 8.710 93.475 8.990 ;
        RECT 93.195 8.310 93.475 8.590 ;
        RECT 95.425 8.710 95.705 8.990 ;
        RECT 95.425 8.310 95.705 8.590 ;
        RECT 78.695 7.125 78.975 7.405 ;
        RECT 79.095 7.125 79.375 7.405 ;
        RECT 79.495 7.125 79.775 7.405 ;
        RECT 192.430 34.960 192.710 35.240 ;
        RECT 192.430 34.560 192.710 34.840 ;
        RECT 192.430 34.160 192.710 34.440 ;
        RECT 199.710 28.050 199.990 28.330 ;
        RECT 199.710 27.650 199.990 27.930 ;
        RECT 199.710 27.250 199.990 27.530 ;
        RECT 200.810 41.415 201.090 41.695 ;
        RECT 200.810 41.015 201.090 41.295 ;
        RECT 200.810 19.030 201.090 19.310 ;
        RECT 200.810 18.630 201.090 18.910 ;
        RECT 200.810 18.230 201.090 18.510 ;
      LAYER met3 ;
        RECT -4.075 108.665 203.595 109.265 ;
        RECT -2.415 107.565 205.835 108.165 ;
        RECT -3.220 97.655 -2.890 98.835 ;
        RECT -4.880 93.980 -4.550 95.160 ;
        RECT -1.290 91.605 -0.690 93.530 ;
        RECT 0.510 80.470 23.110 104.530 ;
        RECT 25.805 80.470 48.405 104.530 ;
        RECT 49.605 80.470 72.205 104.530 ;
        RECT 73.405 80.470 96.005 104.530 ;
        RECT 97.205 80.470 119.805 104.530 ;
        RECT 121.005 80.470 143.605 104.530 ;
        RECT 144.805 80.470 167.405 104.530 ;
        RECT 168.605 91.605 169.205 93.530 ;
        RECT 170.405 80.470 193.005 104.530 ;
        RECT 194.205 91.605 194.805 93.530 ;
        RECT 202.970 85.480 203.570 87.010 ;
        RECT 203.895 85.480 205.835 86.080 ;
        RECT -4.880 78.725 -4.550 79.525 ;
        RECT -4.880 78.395 189.275 78.725 ;
        RECT 133.725 76.425 147.280 77.125 ;
        RECT 133.725 75.880 134.425 76.425 ;
        RECT 168.605 76.240 169.205 76.770 ;
        RECT -2.390 75.010 -1.790 75.410 ;
        RECT 42.690 75.180 134.425 75.880 ;
        RECT 150.090 75.640 189.005 76.240 ;
        RECT -2.390 74.680 0.600 75.010 ;
        RECT 0.930 74.680 42.395 75.010 ;
        RECT 136.120 74.960 189.605 75.290 ;
        RECT 42.690 73.810 130.920 74.510 ;
        RECT 137.595 74.045 189.605 74.375 ;
        RECT 147.920 73.645 148.250 74.045 ;
        RECT 188.175 73.225 188.505 74.045 ;
        RECT 138.580 72.485 138.910 72.905 ;
        RECT 139.440 72.485 139.770 72.905 ;
        RECT 140.300 72.485 140.630 72.905 ;
        RECT 143.830 72.485 144.160 72.905 ;
        RECT 144.690 72.485 145.020 72.905 ;
        RECT 145.550 72.485 145.880 72.885 ;
        RECT -3.220 71.685 -2.890 72.485 ;
        RECT 125.425 72.155 145.880 72.485 ;
        RECT 147.920 71.770 148.250 72.170 ;
        RECT -3.220 71.355 0.605 71.685 ;
        RECT 0.935 71.355 128.475 71.685 ;
        RECT 142.935 71.440 148.250 71.770 ;
        RECT 137.050 70.440 142.080 71.140 ;
        RECT 142.420 70.440 147.370 71.140 ;
        RECT -1.290 69.045 -0.690 69.845 ;
        RECT 194.205 69.045 194.805 69.845 ;
        RECT -1.290 68.715 0.605 69.045 ;
        RECT 0.935 68.715 96.570 69.045 ;
        RECT 124.960 68.715 189.315 69.045 ;
        RECT 189.645 68.715 194.805 69.045 ;
        RECT 0.605 67.785 131.730 68.115 ;
        RECT 189.005 67.915 189.605 68.715 ;
        RECT -4.050 66.705 -3.720 67.505 ;
        RECT 131.995 66.745 147.560 67.445 ;
        RECT -4.050 66.375 0.605 66.705 ;
        RECT 0.935 66.375 131.345 66.705 ;
        RECT 31.700 61.525 32.030 66.375 ;
        RECT 106.370 65.285 110.805 65.615 ;
        RECT 33.400 63.345 144.640 64.045 ;
        RECT 33.400 63.045 38.650 63.345 ;
        RECT 199.550 62.875 200.150 64.000 ;
        RECT 203.895 63.400 205.835 64.000 ;
        RECT 42.650 61.975 144.640 62.675 ;
        RECT 33.665 61.525 34.965 61.535 ;
        RECT 31.700 61.205 34.965 61.525 ;
        RECT 36.995 61.205 38.445 61.535 ;
        RECT 31.700 61.195 33.995 61.205 ;
        RECT 42.650 60.605 144.640 61.305 ;
        RECT 33.400 59.895 38.650 60.195 ;
        RECT 33.400 59.195 40.970 59.895 ;
        RECT 40.270 58.950 40.970 59.195 ;
        RECT 40.270 58.250 46.215 58.950 ;
        RECT 0.605 57.700 1.205 58.230 ;
        RECT 0.605 57.100 188.500 57.700 ;
        RECT 189.005 56.770 189.605 57.300 ;
        RECT 52.850 56.170 189.605 56.770 ;
        RECT 52.850 55.640 53.450 56.170 ;
        RECT 120.535 55.070 186.795 55.670 ;
        RECT 68.215 53.360 79.820 53.690 ;
        RECT 55.800 51.640 118.215 52.640 ;
        RECT 55.800 48.050 95.830 49.050 ;
        RECT 60.410 46.705 60.740 47.105 ;
        RECT 68.090 46.705 68.420 47.105 ;
        RECT 72.650 46.705 72.980 47.105 ;
        RECT 77.210 46.705 77.540 47.105 ;
        RECT 55.415 46.290 58.890 46.620 ;
        RECT 60.410 46.375 77.540 46.705 ;
        RECT 81.770 46.705 82.100 47.105 ;
        RECT 86.330 46.705 86.660 47.105 ;
        RECT 90.890 46.705 91.220 47.105 ;
        RECT 81.770 46.375 91.220 46.705 ;
        RECT 123.190 46.445 132.555 46.775 ;
        RECT 55.415 45.490 55.745 46.290 ;
        RECT 60.435 45.695 84.605 46.025 ;
        RECT 94.015 44.475 118.630 45.475 ;
        RECT 55.800 43.885 93.215 44.385 ;
        RECT 73.115 42.460 100.775 42.790 ;
        RECT 110.690 42.450 111.020 42.850 ;
        RECT 123.190 42.450 123.520 46.445 ;
        RECT 132.225 45.645 132.555 46.445 ;
        RECT 124.280 43.960 144.490 44.960 ;
        RECT 110.690 42.120 125.845 42.450 ;
        RECT 127.875 42.120 129.325 42.450 ;
        RECT 132.225 42.120 136.505 42.450 ;
        RECT 73.120 41.780 100.775 42.110 ;
        RECT 110.690 41.720 111.020 42.120 ;
        RECT 142.835 41.985 189.045 42.585 ;
        RECT 189.645 41.985 191.795 42.585 ;
        RECT 33.875 39.590 35.025 39.970 ;
        RECT 69.010 39.630 90.240 40.630 ;
        RECT 92.215 40.175 118.630 40.675 ;
        RECT 124.280 40.110 144.490 41.110 ;
        RECT 200.650 40.795 201.250 41.920 ;
        RECT 203.895 41.320 205.835 41.920 ;
        RECT 188.175 38.845 188.505 39.665 ;
        RECT 132.560 38.515 188.505 38.845 ;
        RECT 55.440 38.150 95.425 38.480 ;
        RECT 123.495 38.085 130.295 38.415 ;
        RECT 60.435 37.325 71.265 37.655 ;
        RECT 123.495 37.285 123.825 38.085 ;
        RECT 124.125 37.305 127.220 37.635 ;
        RECT 32.775 35.910 33.925 36.290 ;
        RECT 116.215 36.230 129.820 36.965 ;
        RECT 64.575 36.115 129.820 36.230 ;
        RECT 64.575 35.730 118.215 36.115 ;
        RECT 122.365 35.130 122.695 35.530 ;
        RECT 132.560 35.130 132.890 38.515 ;
        RECT 134.940 36.140 144.490 37.140 ;
        RECT 122.365 34.800 126.365 35.130 ;
        RECT 128.075 34.800 136.505 35.130 ;
        RECT 67.610 34.405 91.700 34.735 ;
        RECT 142.835 34.665 189.045 35.265 ;
        RECT 189.645 34.665 192.870 35.265 ;
        RECT 192.270 34.135 192.870 34.665 ;
        RECT 64.575 32.990 118.215 33.490 ;
        RECT 124.730 33.290 129.820 33.740 ;
        RECT 124.730 32.890 144.490 33.290 ;
        RECT -13.115 -45.020 -11.615 32.585 ;
        RECT 53.950 31.745 54.550 32.275 ;
        RECT 80.655 31.950 81.775 32.330 ;
        RECT 128.215 32.290 144.490 32.890 ;
        RECT 128.215 32.165 129.820 32.290 ;
        RECT 52.850 31.145 66.610 31.745 ;
        RECT 124.730 31.315 129.820 32.165 ;
        RECT 92.700 30.765 93.030 31.030 ;
        RECT 120.560 30.765 121.160 31.295 ;
        RECT 52.850 29.645 53.450 30.175 ;
        RECT 92.700 30.165 121.160 30.765 ;
        RECT 124.100 30.645 130.295 30.975 ;
        RECT 92.700 29.900 93.030 30.165 ;
        RECT 52.850 29.045 66.610 29.645 ;
        RECT 124.125 29.585 128.010 29.915 ;
        RECT 129.965 29.845 130.295 30.645 ;
        RECT 80.655 28.460 81.775 28.840 ;
        RECT 124.730 28.395 129.820 29.245 ;
        RECT 134.940 29.200 144.490 30.200 ;
        RECT 199.550 27.825 200.150 28.355 ;
        RECT 64.575 27.300 118.215 27.800 ;
        RECT 124.730 26.820 129.820 27.670 ;
        RECT 131.110 27.360 136.505 27.690 ;
        RECT 67.610 26.055 91.700 26.385 ;
        RECT 123.495 25.760 123.825 26.560 ;
        RECT 123.495 25.430 126.365 25.760 ;
        RECT 128.075 25.430 130.295 25.760 ;
        RECT 64.575 24.560 118.215 25.060 ;
        RECT 116.215 24.445 118.215 24.560 ;
        RECT 116.215 23.595 129.820 24.445 ;
        RECT 132.560 23.610 132.890 27.360 ;
        RECT 142.835 27.225 189.045 27.825 ;
        RECT 189.645 27.225 200.150 27.825 ;
        RECT 134.940 25.350 144.490 26.350 ;
        RECT 60.435 23.135 71.265 23.465 ;
        RECT 132.560 23.280 187.675 23.610 ;
        RECT 123.550 22.925 127.220 23.255 ;
        RECT 55.440 22.310 95.425 22.640 ;
        RECT 69.010 20.160 90.240 21.160 ;
        RECT 92.215 20.115 118.630 20.615 ;
        RECT 73.120 18.680 100.775 19.010 ;
        RECT 110.690 18.670 111.020 19.070 ;
        RECT 123.550 18.670 123.880 22.925 ;
        RECT 128.215 20.180 144.490 21.180 ;
        RECT 200.650 18.805 201.250 19.335 ;
        RECT 110.690 18.340 136.505 18.670 ;
        RECT 73.115 18.000 100.775 18.330 ;
        RECT 110.690 17.940 111.020 18.340 ;
        RECT 142.835 18.205 189.045 18.805 ;
        RECT 189.645 18.205 201.250 18.805 ;
        RECT 55.800 16.405 93.215 16.905 ;
        RECT 134.940 16.330 144.490 17.330 ;
        RECT 94.015 15.315 118.630 16.315 ;
        RECT 55.415 14.500 55.745 15.300 ;
        RECT 60.435 14.765 84.605 15.095 ;
        RECT 55.415 14.170 58.890 14.500 ;
        RECT 60.410 14.085 77.540 14.415 ;
        RECT 60.410 13.685 60.740 14.085 ;
        RECT 68.090 13.685 68.420 14.085 ;
        RECT 72.650 13.685 72.980 14.085 ;
        RECT 77.210 13.685 77.540 14.085 ;
        RECT 81.770 14.085 91.220 14.415 ;
        RECT 81.770 13.685 82.100 14.085 ;
        RECT 86.330 13.685 86.660 14.085 ;
        RECT 90.890 13.685 91.220 14.085 ;
        RECT 55.800 11.740 95.830 12.740 ;
        RECT 55.800 8.150 118.215 9.150 ;
        RECT 68.215 7.100 79.820 7.430 ;
        RECT 35.690 3.500 44.215 6.500 ;
        RECT 47.215 3.500 150.965 6.500 ;
        RECT 35.690 -48.000 38.690 3.500 ;
        RECT 47.215 0.000 143.240 3.000 ;
        RECT 147.965 -48.000 150.965 3.500 ;
      LAYER via3 ;
        RECT 203.905 107.705 204.225 108.025 ;
        RECT 204.305 107.705 204.625 108.025 ;
        RECT 204.705 107.705 205.025 108.025 ;
        RECT 205.105 107.705 205.425 108.025 ;
        RECT 205.505 107.705 205.825 108.025 ;
        RECT -3.215 98.485 -2.895 98.805 ;
        RECT -3.215 98.085 -2.895 98.405 ;
        RECT -3.215 97.685 -2.895 98.005 ;
        RECT -4.875 94.810 -4.555 95.130 ;
        RECT -4.875 94.410 -4.555 94.730 ;
        RECT -4.875 94.010 -4.555 94.330 ;
        RECT -1.150 93.205 -0.830 93.525 ;
        RECT -1.150 92.805 -0.830 93.125 ;
        RECT -1.150 92.405 -0.830 92.725 ;
        RECT -1.150 92.005 -0.830 92.325 ;
        RECT -1.150 91.605 -0.830 91.925 ;
        RECT 0.650 80.570 0.970 80.890 ;
        RECT 1.050 80.570 1.370 80.890 ;
        RECT 1.450 80.570 1.770 80.890 ;
        RECT 1.850 80.570 2.170 80.890 ;
        RECT 2.250 80.570 2.570 80.890 ;
        RECT 2.650 80.570 2.970 80.890 ;
        RECT 3.050 80.570 3.370 80.890 ;
        RECT 3.450 80.570 3.770 80.890 ;
        RECT 3.850 80.570 4.170 80.890 ;
        RECT 4.250 80.570 4.570 80.890 ;
        RECT 4.650 80.570 4.970 80.890 ;
        RECT 5.050 80.570 5.370 80.890 ;
        RECT 5.450 80.570 5.770 80.890 ;
        RECT 5.850 80.570 6.170 80.890 ;
        RECT 6.250 80.570 6.570 80.890 ;
        RECT 6.650 80.570 6.970 80.890 ;
        RECT 7.050 80.570 7.370 80.890 ;
        RECT 7.450 80.570 7.770 80.890 ;
        RECT 7.850 80.570 8.170 80.890 ;
        RECT 8.250 80.570 8.570 80.890 ;
        RECT 8.650 80.570 8.970 80.890 ;
        RECT 9.050 80.570 9.370 80.890 ;
        RECT 9.450 80.570 9.770 80.890 ;
        RECT 9.850 80.570 10.170 80.890 ;
        RECT 10.250 80.570 10.570 80.890 ;
        RECT 10.650 80.570 10.970 80.890 ;
        RECT 11.050 80.570 11.370 80.890 ;
        RECT 11.450 80.570 11.770 80.890 ;
        RECT 11.850 80.570 12.170 80.890 ;
        RECT 12.250 80.570 12.570 80.890 ;
        RECT 12.650 80.570 12.970 80.890 ;
        RECT 13.050 80.570 13.370 80.890 ;
        RECT 13.450 80.570 13.770 80.890 ;
        RECT 13.850 80.570 14.170 80.890 ;
        RECT 14.250 80.570 14.570 80.890 ;
        RECT 14.650 80.570 14.970 80.890 ;
        RECT 15.050 80.570 15.370 80.890 ;
        RECT 15.450 80.570 15.770 80.890 ;
        RECT 15.850 80.570 16.170 80.890 ;
        RECT 16.250 80.570 16.570 80.890 ;
        RECT 16.650 80.570 16.970 80.890 ;
        RECT 17.050 80.570 17.370 80.890 ;
        RECT 17.450 80.570 17.770 80.890 ;
        RECT 17.850 80.570 18.170 80.890 ;
        RECT 18.250 80.570 18.570 80.890 ;
        RECT 18.650 80.570 18.970 80.890 ;
        RECT 19.050 80.570 19.370 80.890 ;
        RECT 19.450 80.570 19.770 80.890 ;
        RECT 19.850 80.570 20.170 80.890 ;
        RECT 20.250 80.570 20.570 80.890 ;
        RECT 20.650 80.570 20.970 80.890 ;
        RECT 21.050 80.570 21.370 80.890 ;
        RECT 21.450 80.570 21.770 80.890 ;
        RECT 21.850 80.570 22.170 80.890 ;
        RECT 22.250 80.570 22.570 80.890 ;
        RECT 22.650 80.570 22.970 80.890 ;
        RECT 25.945 80.570 26.265 80.890 ;
        RECT 26.345 80.570 26.665 80.890 ;
        RECT 26.745 80.570 27.065 80.890 ;
        RECT 27.145 80.570 27.465 80.890 ;
        RECT 27.545 80.570 27.865 80.890 ;
        RECT 27.945 80.570 28.265 80.890 ;
        RECT 28.345 80.570 28.665 80.890 ;
        RECT 28.745 80.570 29.065 80.890 ;
        RECT 29.145 80.570 29.465 80.890 ;
        RECT 29.545 80.570 29.865 80.890 ;
        RECT 29.945 80.570 30.265 80.890 ;
        RECT 30.345 80.570 30.665 80.890 ;
        RECT 30.745 80.570 31.065 80.890 ;
        RECT 31.145 80.570 31.465 80.890 ;
        RECT 31.545 80.570 31.865 80.890 ;
        RECT 31.945 80.570 32.265 80.890 ;
        RECT 32.345 80.570 32.665 80.890 ;
        RECT 32.745 80.570 33.065 80.890 ;
        RECT 33.145 80.570 33.465 80.890 ;
        RECT 33.545 80.570 33.865 80.890 ;
        RECT 33.945 80.570 34.265 80.890 ;
        RECT 34.345 80.570 34.665 80.890 ;
        RECT 34.745 80.570 35.065 80.890 ;
        RECT 35.145 80.570 35.465 80.890 ;
        RECT 35.545 80.570 35.865 80.890 ;
        RECT 35.945 80.570 36.265 80.890 ;
        RECT 36.345 80.570 36.665 80.890 ;
        RECT 36.745 80.570 37.065 80.890 ;
        RECT 37.145 80.570 37.465 80.890 ;
        RECT 37.545 80.570 37.865 80.890 ;
        RECT 37.945 80.570 38.265 80.890 ;
        RECT 38.345 80.570 38.665 80.890 ;
        RECT 38.745 80.570 39.065 80.890 ;
        RECT 39.145 80.570 39.465 80.890 ;
        RECT 39.545 80.570 39.865 80.890 ;
        RECT 39.945 80.570 40.265 80.890 ;
        RECT 40.345 80.570 40.665 80.890 ;
        RECT 40.745 80.570 41.065 80.890 ;
        RECT 41.145 80.570 41.465 80.890 ;
        RECT 41.545 80.570 41.865 80.890 ;
        RECT 41.945 80.570 42.265 80.890 ;
        RECT 42.345 80.570 42.665 80.890 ;
        RECT 42.745 80.570 43.065 80.890 ;
        RECT 43.145 80.570 43.465 80.890 ;
        RECT 43.545 80.570 43.865 80.890 ;
        RECT 43.945 80.570 44.265 80.890 ;
        RECT 44.345 80.570 44.665 80.890 ;
        RECT 44.745 80.570 45.065 80.890 ;
        RECT 45.145 80.570 45.465 80.890 ;
        RECT 45.545 80.570 45.865 80.890 ;
        RECT 45.945 80.570 46.265 80.890 ;
        RECT 46.345 80.570 46.665 80.890 ;
        RECT 46.745 80.570 47.065 80.890 ;
        RECT 47.145 80.570 47.465 80.890 ;
        RECT 47.545 80.570 47.865 80.890 ;
        RECT 47.945 80.570 48.265 80.890 ;
        RECT 49.745 80.570 50.065 80.890 ;
        RECT 50.145 80.570 50.465 80.890 ;
        RECT 50.545 80.570 50.865 80.890 ;
        RECT 50.945 80.570 51.265 80.890 ;
        RECT 51.345 80.570 51.665 80.890 ;
        RECT 51.745 80.570 52.065 80.890 ;
        RECT 52.145 80.570 52.465 80.890 ;
        RECT 52.545 80.570 52.865 80.890 ;
        RECT 52.945 80.570 53.265 80.890 ;
        RECT 53.345 80.570 53.665 80.890 ;
        RECT 53.745 80.570 54.065 80.890 ;
        RECT 54.145 80.570 54.465 80.890 ;
        RECT 54.545 80.570 54.865 80.890 ;
        RECT 54.945 80.570 55.265 80.890 ;
        RECT 55.345 80.570 55.665 80.890 ;
        RECT 55.745 80.570 56.065 80.890 ;
        RECT 56.145 80.570 56.465 80.890 ;
        RECT 56.545 80.570 56.865 80.890 ;
        RECT 56.945 80.570 57.265 80.890 ;
        RECT 57.345 80.570 57.665 80.890 ;
        RECT 57.745 80.570 58.065 80.890 ;
        RECT 58.145 80.570 58.465 80.890 ;
        RECT 58.545 80.570 58.865 80.890 ;
        RECT 58.945 80.570 59.265 80.890 ;
        RECT 59.345 80.570 59.665 80.890 ;
        RECT 59.745 80.570 60.065 80.890 ;
        RECT 60.145 80.570 60.465 80.890 ;
        RECT 60.545 80.570 60.865 80.890 ;
        RECT 60.945 80.570 61.265 80.890 ;
        RECT 61.345 80.570 61.665 80.890 ;
        RECT 61.745 80.570 62.065 80.890 ;
        RECT 62.145 80.570 62.465 80.890 ;
        RECT 62.545 80.570 62.865 80.890 ;
        RECT 62.945 80.570 63.265 80.890 ;
        RECT 63.345 80.570 63.665 80.890 ;
        RECT 63.745 80.570 64.065 80.890 ;
        RECT 64.145 80.570 64.465 80.890 ;
        RECT 64.545 80.570 64.865 80.890 ;
        RECT 64.945 80.570 65.265 80.890 ;
        RECT 65.345 80.570 65.665 80.890 ;
        RECT 65.745 80.570 66.065 80.890 ;
        RECT 66.145 80.570 66.465 80.890 ;
        RECT 66.545 80.570 66.865 80.890 ;
        RECT 66.945 80.570 67.265 80.890 ;
        RECT 67.345 80.570 67.665 80.890 ;
        RECT 67.745 80.570 68.065 80.890 ;
        RECT 68.145 80.570 68.465 80.890 ;
        RECT 68.545 80.570 68.865 80.890 ;
        RECT 68.945 80.570 69.265 80.890 ;
        RECT 69.345 80.570 69.665 80.890 ;
        RECT 69.745 80.570 70.065 80.890 ;
        RECT 70.145 80.570 70.465 80.890 ;
        RECT 70.545 80.570 70.865 80.890 ;
        RECT 70.945 80.570 71.265 80.890 ;
        RECT 71.345 80.570 71.665 80.890 ;
        RECT 71.745 80.570 72.065 80.890 ;
        RECT 73.545 80.570 73.865 80.890 ;
        RECT 73.945 80.570 74.265 80.890 ;
        RECT 74.345 80.570 74.665 80.890 ;
        RECT 74.745 80.570 75.065 80.890 ;
        RECT 75.145 80.570 75.465 80.890 ;
        RECT 75.545 80.570 75.865 80.890 ;
        RECT 75.945 80.570 76.265 80.890 ;
        RECT 76.345 80.570 76.665 80.890 ;
        RECT 76.745 80.570 77.065 80.890 ;
        RECT 77.145 80.570 77.465 80.890 ;
        RECT 77.545 80.570 77.865 80.890 ;
        RECT 77.945 80.570 78.265 80.890 ;
        RECT 78.345 80.570 78.665 80.890 ;
        RECT 78.745 80.570 79.065 80.890 ;
        RECT 79.145 80.570 79.465 80.890 ;
        RECT 79.545 80.570 79.865 80.890 ;
        RECT 79.945 80.570 80.265 80.890 ;
        RECT 80.345 80.570 80.665 80.890 ;
        RECT 80.745 80.570 81.065 80.890 ;
        RECT 81.145 80.570 81.465 80.890 ;
        RECT 81.545 80.570 81.865 80.890 ;
        RECT 81.945 80.570 82.265 80.890 ;
        RECT 82.345 80.570 82.665 80.890 ;
        RECT 82.745 80.570 83.065 80.890 ;
        RECT 83.145 80.570 83.465 80.890 ;
        RECT 83.545 80.570 83.865 80.890 ;
        RECT 83.945 80.570 84.265 80.890 ;
        RECT 84.345 80.570 84.665 80.890 ;
        RECT 84.745 80.570 85.065 80.890 ;
        RECT 85.145 80.570 85.465 80.890 ;
        RECT 85.545 80.570 85.865 80.890 ;
        RECT 85.945 80.570 86.265 80.890 ;
        RECT 86.345 80.570 86.665 80.890 ;
        RECT 86.745 80.570 87.065 80.890 ;
        RECT 87.145 80.570 87.465 80.890 ;
        RECT 87.545 80.570 87.865 80.890 ;
        RECT 87.945 80.570 88.265 80.890 ;
        RECT 88.345 80.570 88.665 80.890 ;
        RECT 88.745 80.570 89.065 80.890 ;
        RECT 89.145 80.570 89.465 80.890 ;
        RECT 89.545 80.570 89.865 80.890 ;
        RECT 89.945 80.570 90.265 80.890 ;
        RECT 90.345 80.570 90.665 80.890 ;
        RECT 90.745 80.570 91.065 80.890 ;
        RECT 91.145 80.570 91.465 80.890 ;
        RECT 91.545 80.570 91.865 80.890 ;
        RECT 91.945 80.570 92.265 80.890 ;
        RECT 92.345 80.570 92.665 80.890 ;
        RECT 92.745 80.570 93.065 80.890 ;
        RECT 93.145 80.570 93.465 80.890 ;
        RECT 93.545 80.570 93.865 80.890 ;
        RECT 93.945 80.570 94.265 80.890 ;
        RECT 94.345 80.570 94.665 80.890 ;
        RECT 94.745 80.570 95.065 80.890 ;
        RECT 95.145 80.570 95.465 80.890 ;
        RECT 95.545 80.570 95.865 80.890 ;
        RECT 97.345 80.570 97.665 80.890 ;
        RECT 97.745 80.570 98.065 80.890 ;
        RECT 98.145 80.570 98.465 80.890 ;
        RECT 98.545 80.570 98.865 80.890 ;
        RECT 98.945 80.570 99.265 80.890 ;
        RECT 99.345 80.570 99.665 80.890 ;
        RECT 99.745 80.570 100.065 80.890 ;
        RECT 100.145 80.570 100.465 80.890 ;
        RECT 100.545 80.570 100.865 80.890 ;
        RECT 100.945 80.570 101.265 80.890 ;
        RECT 101.345 80.570 101.665 80.890 ;
        RECT 101.745 80.570 102.065 80.890 ;
        RECT 102.145 80.570 102.465 80.890 ;
        RECT 102.545 80.570 102.865 80.890 ;
        RECT 102.945 80.570 103.265 80.890 ;
        RECT 103.345 80.570 103.665 80.890 ;
        RECT 103.745 80.570 104.065 80.890 ;
        RECT 104.145 80.570 104.465 80.890 ;
        RECT 104.545 80.570 104.865 80.890 ;
        RECT 104.945 80.570 105.265 80.890 ;
        RECT 105.345 80.570 105.665 80.890 ;
        RECT 105.745 80.570 106.065 80.890 ;
        RECT 106.145 80.570 106.465 80.890 ;
        RECT 106.545 80.570 106.865 80.890 ;
        RECT 106.945 80.570 107.265 80.890 ;
        RECT 107.345 80.570 107.665 80.890 ;
        RECT 107.745 80.570 108.065 80.890 ;
        RECT 108.145 80.570 108.465 80.890 ;
        RECT 108.545 80.570 108.865 80.890 ;
        RECT 108.945 80.570 109.265 80.890 ;
        RECT 109.345 80.570 109.665 80.890 ;
        RECT 109.745 80.570 110.065 80.890 ;
        RECT 110.145 80.570 110.465 80.890 ;
        RECT 110.545 80.570 110.865 80.890 ;
        RECT 110.945 80.570 111.265 80.890 ;
        RECT 111.345 80.570 111.665 80.890 ;
        RECT 111.745 80.570 112.065 80.890 ;
        RECT 112.145 80.570 112.465 80.890 ;
        RECT 112.545 80.570 112.865 80.890 ;
        RECT 112.945 80.570 113.265 80.890 ;
        RECT 113.345 80.570 113.665 80.890 ;
        RECT 113.745 80.570 114.065 80.890 ;
        RECT 114.145 80.570 114.465 80.890 ;
        RECT 114.545 80.570 114.865 80.890 ;
        RECT 114.945 80.570 115.265 80.890 ;
        RECT 115.345 80.570 115.665 80.890 ;
        RECT 115.745 80.570 116.065 80.890 ;
        RECT 116.145 80.570 116.465 80.890 ;
        RECT 116.545 80.570 116.865 80.890 ;
        RECT 116.945 80.570 117.265 80.890 ;
        RECT 117.345 80.570 117.665 80.890 ;
        RECT 117.745 80.570 118.065 80.890 ;
        RECT 118.145 80.570 118.465 80.890 ;
        RECT 118.545 80.570 118.865 80.890 ;
        RECT 118.945 80.570 119.265 80.890 ;
        RECT 119.345 80.570 119.665 80.890 ;
        RECT 121.145 80.570 121.465 80.890 ;
        RECT 121.545 80.570 121.865 80.890 ;
        RECT 121.945 80.570 122.265 80.890 ;
        RECT 122.345 80.570 122.665 80.890 ;
        RECT 122.745 80.570 123.065 80.890 ;
        RECT 123.145 80.570 123.465 80.890 ;
        RECT 123.545 80.570 123.865 80.890 ;
        RECT 123.945 80.570 124.265 80.890 ;
        RECT 124.345 80.570 124.665 80.890 ;
        RECT 124.745 80.570 125.065 80.890 ;
        RECT 125.145 80.570 125.465 80.890 ;
        RECT 125.545 80.570 125.865 80.890 ;
        RECT 125.945 80.570 126.265 80.890 ;
        RECT 126.345 80.570 126.665 80.890 ;
        RECT 126.745 80.570 127.065 80.890 ;
        RECT 127.145 80.570 127.465 80.890 ;
        RECT 127.545 80.570 127.865 80.890 ;
        RECT 127.945 80.570 128.265 80.890 ;
        RECT 128.345 80.570 128.665 80.890 ;
        RECT 128.745 80.570 129.065 80.890 ;
        RECT 129.145 80.570 129.465 80.890 ;
        RECT 129.545 80.570 129.865 80.890 ;
        RECT 129.945 80.570 130.265 80.890 ;
        RECT 130.345 80.570 130.665 80.890 ;
        RECT 130.745 80.570 131.065 80.890 ;
        RECT 131.145 80.570 131.465 80.890 ;
        RECT 131.545 80.570 131.865 80.890 ;
        RECT 131.945 80.570 132.265 80.890 ;
        RECT 132.345 80.570 132.665 80.890 ;
        RECT 132.745 80.570 133.065 80.890 ;
        RECT 133.145 80.570 133.465 80.890 ;
        RECT 133.545 80.570 133.865 80.890 ;
        RECT 133.945 80.570 134.265 80.890 ;
        RECT 134.345 80.570 134.665 80.890 ;
        RECT 134.745 80.570 135.065 80.890 ;
        RECT 135.145 80.570 135.465 80.890 ;
        RECT 135.545 80.570 135.865 80.890 ;
        RECT 135.945 80.570 136.265 80.890 ;
        RECT 136.345 80.570 136.665 80.890 ;
        RECT 136.745 80.570 137.065 80.890 ;
        RECT 137.145 80.570 137.465 80.890 ;
        RECT 137.545 80.570 137.865 80.890 ;
        RECT 137.945 80.570 138.265 80.890 ;
        RECT 138.345 80.570 138.665 80.890 ;
        RECT 138.745 80.570 139.065 80.890 ;
        RECT 139.145 80.570 139.465 80.890 ;
        RECT 139.545 80.570 139.865 80.890 ;
        RECT 139.945 80.570 140.265 80.890 ;
        RECT 140.345 80.570 140.665 80.890 ;
        RECT 140.745 80.570 141.065 80.890 ;
        RECT 141.145 80.570 141.465 80.890 ;
        RECT 141.545 80.570 141.865 80.890 ;
        RECT 141.945 80.570 142.265 80.890 ;
        RECT 142.345 80.570 142.665 80.890 ;
        RECT 142.745 80.570 143.065 80.890 ;
        RECT 143.145 80.570 143.465 80.890 ;
        RECT 168.745 93.205 169.065 93.525 ;
        RECT 168.745 92.805 169.065 93.125 ;
        RECT 168.745 92.405 169.065 92.725 ;
        RECT 168.745 92.005 169.065 92.325 ;
        RECT 168.745 91.605 169.065 91.925 ;
        RECT 144.945 80.570 145.265 80.890 ;
        RECT 145.345 80.570 145.665 80.890 ;
        RECT 145.745 80.570 146.065 80.890 ;
        RECT 146.145 80.570 146.465 80.890 ;
        RECT 146.545 80.570 146.865 80.890 ;
        RECT 146.945 80.570 147.265 80.890 ;
        RECT 147.345 80.570 147.665 80.890 ;
        RECT 147.745 80.570 148.065 80.890 ;
        RECT 148.145 80.570 148.465 80.890 ;
        RECT 148.545 80.570 148.865 80.890 ;
        RECT 148.945 80.570 149.265 80.890 ;
        RECT 149.345 80.570 149.665 80.890 ;
        RECT 149.745 80.570 150.065 80.890 ;
        RECT 150.145 80.570 150.465 80.890 ;
        RECT 150.545 80.570 150.865 80.890 ;
        RECT 150.945 80.570 151.265 80.890 ;
        RECT 151.345 80.570 151.665 80.890 ;
        RECT 151.745 80.570 152.065 80.890 ;
        RECT 152.145 80.570 152.465 80.890 ;
        RECT 152.545 80.570 152.865 80.890 ;
        RECT 152.945 80.570 153.265 80.890 ;
        RECT 153.345 80.570 153.665 80.890 ;
        RECT 153.745 80.570 154.065 80.890 ;
        RECT 154.145 80.570 154.465 80.890 ;
        RECT 154.545 80.570 154.865 80.890 ;
        RECT 154.945 80.570 155.265 80.890 ;
        RECT 155.345 80.570 155.665 80.890 ;
        RECT 155.745 80.570 156.065 80.890 ;
        RECT 156.145 80.570 156.465 80.890 ;
        RECT 156.545 80.570 156.865 80.890 ;
        RECT 156.945 80.570 157.265 80.890 ;
        RECT 157.345 80.570 157.665 80.890 ;
        RECT 157.745 80.570 158.065 80.890 ;
        RECT 158.145 80.570 158.465 80.890 ;
        RECT 158.545 80.570 158.865 80.890 ;
        RECT 158.945 80.570 159.265 80.890 ;
        RECT 159.345 80.570 159.665 80.890 ;
        RECT 159.745 80.570 160.065 80.890 ;
        RECT 160.145 80.570 160.465 80.890 ;
        RECT 160.545 80.570 160.865 80.890 ;
        RECT 160.945 80.570 161.265 80.890 ;
        RECT 161.345 80.570 161.665 80.890 ;
        RECT 161.745 80.570 162.065 80.890 ;
        RECT 162.145 80.570 162.465 80.890 ;
        RECT 162.545 80.570 162.865 80.890 ;
        RECT 162.945 80.570 163.265 80.890 ;
        RECT 163.345 80.570 163.665 80.890 ;
        RECT 163.745 80.570 164.065 80.890 ;
        RECT 164.145 80.570 164.465 80.890 ;
        RECT 164.545 80.570 164.865 80.890 ;
        RECT 164.945 80.570 165.265 80.890 ;
        RECT 165.345 80.570 165.665 80.890 ;
        RECT 165.745 80.570 166.065 80.890 ;
        RECT 166.145 80.570 166.465 80.890 ;
        RECT 166.545 80.570 166.865 80.890 ;
        RECT 166.945 80.570 167.265 80.890 ;
        RECT 194.345 93.205 194.665 93.525 ;
        RECT 194.345 92.805 194.665 93.125 ;
        RECT 194.345 92.405 194.665 92.725 ;
        RECT 194.345 92.005 194.665 92.325 ;
        RECT 194.345 91.605 194.665 91.925 ;
        RECT 203.110 86.685 203.430 87.005 ;
        RECT 203.110 86.285 203.430 86.605 ;
        RECT 203.110 85.885 203.430 86.205 ;
        RECT 203.110 85.485 203.430 85.805 ;
        RECT 203.905 85.620 204.225 85.940 ;
        RECT 204.305 85.620 204.625 85.940 ;
        RECT 204.705 85.620 205.025 85.940 ;
        RECT 205.105 85.620 205.425 85.940 ;
        RECT 205.505 85.620 205.825 85.940 ;
        RECT 170.545 80.570 170.865 80.890 ;
        RECT 170.945 80.570 171.265 80.890 ;
        RECT 171.345 80.570 171.665 80.890 ;
        RECT 171.745 80.570 172.065 80.890 ;
        RECT 172.145 80.570 172.465 80.890 ;
        RECT 172.545 80.570 172.865 80.890 ;
        RECT 172.945 80.570 173.265 80.890 ;
        RECT 173.345 80.570 173.665 80.890 ;
        RECT 173.745 80.570 174.065 80.890 ;
        RECT 174.145 80.570 174.465 80.890 ;
        RECT 174.545 80.570 174.865 80.890 ;
        RECT 174.945 80.570 175.265 80.890 ;
        RECT 175.345 80.570 175.665 80.890 ;
        RECT 175.745 80.570 176.065 80.890 ;
        RECT 176.145 80.570 176.465 80.890 ;
        RECT 176.545 80.570 176.865 80.890 ;
        RECT 176.945 80.570 177.265 80.890 ;
        RECT 177.345 80.570 177.665 80.890 ;
        RECT 177.745 80.570 178.065 80.890 ;
        RECT 178.145 80.570 178.465 80.890 ;
        RECT 178.545 80.570 178.865 80.890 ;
        RECT 178.945 80.570 179.265 80.890 ;
        RECT 179.345 80.570 179.665 80.890 ;
        RECT 179.745 80.570 180.065 80.890 ;
        RECT 180.145 80.570 180.465 80.890 ;
        RECT 180.545 80.570 180.865 80.890 ;
        RECT 180.945 80.570 181.265 80.890 ;
        RECT 181.345 80.570 181.665 80.890 ;
        RECT 181.745 80.570 182.065 80.890 ;
        RECT 182.145 80.570 182.465 80.890 ;
        RECT 182.545 80.570 182.865 80.890 ;
        RECT 182.945 80.570 183.265 80.890 ;
        RECT 183.345 80.570 183.665 80.890 ;
        RECT 183.745 80.570 184.065 80.890 ;
        RECT 184.145 80.570 184.465 80.890 ;
        RECT 184.545 80.570 184.865 80.890 ;
        RECT 184.945 80.570 185.265 80.890 ;
        RECT 185.345 80.570 185.665 80.890 ;
        RECT 185.745 80.570 186.065 80.890 ;
        RECT 186.145 80.570 186.465 80.890 ;
        RECT 186.545 80.570 186.865 80.890 ;
        RECT 186.945 80.570 187.265 80.890 ;
        RECT 187.345 80.570 187.665 80.890 ;
        RECT 187.745 80.570 188.065 80.890 ;
        RECT 188.145 80.570 188.465 80.890 ;
        RECT 188.545 80.570 188.865 80.890 ;
        RECT 188.945 80.570 189.265 80.890 ;
        RECT 189.345 80.570 189.665 80.890 ;
        RECT 189.745 80.570 190.065 80.890 ;
        RECT 190.145 80.570 190.465 80.890 ;
        RECT 190.545 80.570 190.865 80.890 ;
        RECT 190.945 80.570 191.265 80.890 ;
        RECT 191.345 80.570 191.665 80.890 ;
        RECT 191.745 80.570 192.065 80.890 ;
        RECT 192.145 80.570 192.465 80.890 ;
        RECT 192.545 80.570 192.865 80.890 ;
        RECT 140.255 76.615 140.575 76.935 ;
        RECT 140.655 76.615 140.975 76.935 ;
        RECT 141.055 76.615 141.375 76.935 ;
        RECT 141.455 76.615 141.775 76.935 ;
        RECT 141.855 76.615 142.175 76.935 ;
        RECT 44.255 75.370 44.575 75.690 ;
        RECT 44.655 75.370 44.975 75.690 ;
        RECT 45.055 75.370 45.375 75.690 ;
        RECT 45.455 75.370 45.775 75.690 ;
        RECT 45.855 75.370 46.175 75.690 ;
        RECT 68.255 75.370 68.575 75.690 ;
        RECT 68.655 75.370 68.975 75.690 ;
        RECT 69.055 75.370 69.375 75.690 ;
        RECT 69.455 75.370 69.775 75.690 ;
        RECT 69.855 75.370 70.175 75.690 ;
        RECT 92.255 75.370 92.575 75.690 ;
        RECT 92.655 75.370 92.975 75.690 ;
        RECT 93.055 75.370 93.375 75.690 ;
        RECT 93.455 75.370 93.775 75.690 ;
        RECT 93.855 75.370 94.175 75.690 ;
        RECT 116.255 75.370 116.575 75.690 ;
        RECT 116.655 75.370 116.975 75.690 ;
        RECT 117.055 75.370 117.375 75.690 ;
        RECT 117.455 75.370 117.775 75.690 ;
        RECT 117.855 75.370 118.175 75.690 ;
        RECT 44.255 74.000 44.575 74.320 ;
        RECT 44.655 74.000 44.975 74.320 ;
        RECT 45.055 74.000 45.375 74.320 ;
        RECT 45.455 74.000 45.775 74.320 ;
        RECT 45.855 74.000 46.175 74.320 ;
        RECT 68.255 74.000 68.575 74.320 ;
        RECT 68.655 74.000 68.975 74.320 ;
        RECT 69.055 74.000 69.375 74.320 ;
        RECT 69.455 74.000 69.775 74.320 ;
        RECT 69.855 74.000 70.175 74.320 ;
        RECT 92.255 74.000 92.575 74.320 ;
        RECT 92.655 74.000 92.975 74.320 ;
        RECT 93.055 74.000 93.375 74.320 ;
        RECT 93.455 74.000 93.775 74.320 ;
        RECT 93.855 74.000 94.175 74.320 ;
        RECT 116.255 74.000 116.575 74.320 ;
        RECT 116.655 74.000 116.975 74.320 ;
        RECT 117.055 74.000 117.375 74.320 ;
        RECT 117.455 74.000 117.775 74.320 ;
        RECT 117.855 74.000 118.175 74.320 ;
        RECT 56.255 63.535 56.575 63.855 ;
        RECT 56.655 63.535 56.975 63.855 ;
        RECT 57.055 63.535 57.375 63.855 ;
        RECT 57.455 63.535 57.775 63.855 ;
        RECT 57.855 63.535 58.175 63.855 ;
        RECT 80.255 63.535 80.575 63.855 ;
        RECT 80.655 63.535 80.975 63.855 ;
        RECT 81.055 63.535 81.375 63.855 ;
        RECT 81.455 63.535 81.775 63.855 ;
        RECT 81.855 63.535 82.175 63.855 ;
        RECT 104.255 63.535 104.575 63.855 ;
        RECT 104.655 63.535 104.975 63.855 ;
        RECT 105.055 63.535 105.375 63.855 ;
        RECT 105.455 63.535 105.775 63.855 ;
        RECT 105.855 63.535 106.175 63.855 ;
        RECT 128.255 63.535 128.575 63.855 ;
        RECT 128.655 63.535 128.975 63.855 ;
        RECT 129.055 63.535 129.375 63.855 ;
        RECT 129.455 63.535 129.775 63.855 ;
        RECT 129.855 63.535 130.175 63.855 ;
        RECT 199.690 63.675 200.010 63.995 ;
        RECT 199.690 63.275 200.010 63.595 ;
        RECT 203.905 63.540 204.225 63.860 ;
        RECT 204.305 63.540 204.625 63.860 ;
        RECT 204.705 63.540 205.025 63.860 ;
        RECT 205.105 63.540 205.425 63.860 ;
        RECT 205.505 63.540 205.825 63.860 ;
        RECT 199.690 62.875 200.010 63.195 ;
        RECT 56.255 62.165 56.575 62.485 ;
        RECT 56.655 62.165 56.975 62.485 ;
        RECT 57.055 62.165 57.375 62.485 ;
        RECT 57.455 62.165 57.775 62.485 ;
        RECT 57.855 62.165 58.175 62.485 ;
        RECT 80.255 62.165 80.575 62.485 ;
        RECT 80.655 62.165 80.975 62.485 ;
        RECT 81.055 62.165 81.375 62.485 ;
        RECT 81.455 62.165 81.775 62.485 ;
        RECT 81.855 62.165 82.175 62.485 ;
        RECT 104.255 62.165 104.575 62.485 ;
        RECT 104.655 62.165 104.975 62.485 ;
        RECT 105.055 62.165 105.375 62.485 ;
        RECT 105.455 62.165 105.775 62.485 ;
        RECT 105.855 62.165 106.175 62.485 ;
        RECT 128.255 62.165 128.575 62.485 ;
        RECT 128.655 62.165 128.975 62.485 ;
        RECT 129.055 62.165 129.375 62.485 ;
        RECT 129.455 62.165 129.775 62.485 ;
        RECT 129.855 62.165 130.175 62.485 ;
        RECT 56.255 60.795 56.575 61.115 ;
        RECT 56.655 60.795 56.975 61.115 ;
        RECT 57.055 60.795 57.375 61.115 ;
        RECT 57.455 60.795 57.775 61.115 ;
        RECT 57.855 60.795 58.175 61.115 ;
        RECT 80.255 60.795 80.575 61.115 ;
        RECT 80.655 60.795 80.975 61.115 ;
        RECT 81.055 60.795 81.375 61.115 ;
        RECT 81.455 60.795 81.775 61.115 ;
        RECT 81.855 60.795 82.175 61.115 ;
        RECT 104.255 60.795 104.575 61.115 ;
        RECT 104.655 60.795 104.975 61.115 ;
        RECT 105.055 60.795 105.375 61.115 ;
        RECT 105.455 60.795 105.775 61.115 ;
        RECT 105.855 60.795 106.175 61.115 ;
        RECT 128.255 60.795 128.575 61.115 ;
        RECT 128.655 60.795 128.975 61.115 ;
        RECT 129.055 60.795 129.375 61.115 ;
        RECT 129.455 60.795 129.775 61.115 ;
        RECT 129.855 60.795 130.175 61.115 ;
        RECT 44.255 58.440 44.575 58.760 ;
        RECT 44.655 58.440 44.975 58.760 ;
        RECT 45.055 58.440 45.375 58.760 ;
        RECT 45.455 58.440 45.775 58.760 ;
        RECT 45.855 58.440 46.175 58.760 ;
        RECT 68.655 53.365 68.975 53.685 ;
        RECT 69.055 53.365 69.375 53.685 ;
        RECT 69.455 53.365 69.775 53.685 ;
        RECT 56.255 51.780 58.175 52.500 ;
        RECT 80.255 51.780 82.175 52.500 ;
        RECT 104.255 51.780 106.175 52.500 ;
        RECT 56.255 48.190 58.175 48.910 ;
        RECT 80.255 48.190 82.175 48.910 ;
        RECT 104.255 44.615 106.175 45.335 ;
        RECT 68.255 43.975 68.575 44.295 ;
        RECT 68.655 43.975 68.975 44.295 ;
        RECT 69.055 43.975 69.375 44.295 ;
        RECT 69.455 43.975 69.775 44.295 ;
        RECT 69.855 43.975 70.175 44.295 ;
        RECT 92.255 43.975 92.575 44.295 ;
        RECT 92.655 43.975 92.975 44.295 ;
        RECT 128.255 44.100 130.175 44.820 ;
        RECT 200.790 41.595 201.110 41.915 ;
        RECT 200.790 41.195 201.110 41.515 ;
        RECT 203.905 41.460 204.225 41.780 ;
        RECT 204.305 41.460 204.625 41.780 ;
        RECT 204.705 41.460 205.025 41.780 ;
        RECT 205.105 41.460 205.425 41.780 ;
        RECT 205.505 41.460 205.825 41.780 ;
        RECT 33.905 39.620 34.225 39.940 ;
        RECT 34.305 39.620 34.625 39.940 ;
        RECT 34.705 39.620 35.025 39.940 ;
        RECT 80.255 39.770 82.175 40.490 ;
        RECT 92.255 40.265 92.575 40.585 ;
        RECT 92.655 40.265 92.975 40.585 ;
        RECT 93.055 40.265 93.375 40.585 ;
        RECT 93.455 40.265 93.775 40.585 ;
        RECT 93.855 40.265 94.175 40.585 ;
        RECT 116.255 40.265 116.575 40.585 ;
        RECT 116.655 40.265 116.975 40.585 ;
        RECT 117.055 40.265 117.375 40.585 ;
        RECT 117.455 40.265 117.775 40.585 ;
        RECT 117.855 40.265 118.175 40.585 ;
        RECT 140.255 40.250 142.175 40.970 ;
        RECT 200.790 40.795 201.110 41.115 ;
        RECT 116.255 36.460 116.575 36.780 ;
        RECT 116.655 36.460 116.975 36.780 ;
        RECT 117.055 36.460 117.375 36.780 ;
        RECT 117.455 36.460 117.775 36.780 ;
        RECT 117.855 36.460 118.175 36.780 ;
        RECT 32.805 35.940 33.125 36.260 ;
        RECT 33.205 35.940 33.525 36.260 ;
        RECT 33.605 35.940 33.925 36.260 ;
        RECT 124.930 36.180 125.650 36.900 ;
        RECT 68.255 35.820 68.575 36.140 ;
        RECT 68.655 35.820 68.975 36.140 ;
        RECT 69.055 35.820 69.375 36.140 ;
        RECT 69.455 35.820 69.775 36.140 ;
        RECT 69.855 35.820 70.175 36.140 ;
        RECT 92.255 35.820 92.575 36.140 ;
        RECT 92.655 35.820 92.975 36.140 ;
        RECT 93.055 35.820 93.375 36.140 ;
        RECT 93.455 35.820 93.775 36.140 ;
        RECT 93.855 35.820 94.175 36.140 ;
        RECT 116.255 35.820 116.575 36.140 ;
        RECT 116.655 35.820 116.975 36.140 ;
        RECT 117.055 35.820 117.375 36.140 ;
        RECT 117.455 35.820 117.775 36.140 ;
        RECT 117.855 35.820 118.175 36.140 ;
        RECT 140.255 36.280 142.175 37.000 ;
        RECT 68.255 33.080 68.575 33.400 ;
        RECT 68.655 33.080 68.975 33.400 ;
        RECT 69.055 33.080 69.375 33.400 ;
        RECT 69.455 33.080 69.775 33.400 ;
        RECT 69.855 33.080 70.175 33.400 ;
        RECT 92.255 33.080 92.575 33.400 ;
        RECT 92.655 33.080 92.975 33.400 ;
        RECT 93.055 33.080 93.375 33.400 ;
        RECT 93.455 33.080 93.775 33.400 ;
        RECT 93.855 33.080 94.175 33.400 ;
        RECT 116.255 33.080 116.575 33.400 ;
        RECT 116.655 33.080 116.975 33.400 ;
        RECT 117.055 33.080 117.375 33.400 ;
        RECT 117.455 33.080 117.775 33.400 ;
        RECT 117.855 33.080 118.175 33.400 ;
        RECT 128.930 32.955 129.650 33.675 ;
        RECT -12.925 32.260 -12.605 32.580 ;
        RECT -12.525 32.260 -12.205 32.580 ;
        RECT -12.125 32.260 -11.805 32.580 ;
        RECT 80.655 31.980 80.975 32.300 ;
        RECT 81.055 31.980 81.375 32.300 ;
        RECT 81.455 31.980 81.775 32.300 ;
        RECT 128.930 31.380 129.650 32.100 ;
        RECT -12.925 28.580 -12.605 28.900 ;
        RECT -12.525 28.580 -12.205 28.900 ;
        RECT -12.125 28.580 -11.805 28.900 ;
        RECT 80.655 28.490 80.975 28.810 ;
        RECT 81.055 28.490 81.375 28.810 ;
        RECT 81.455 28.490 81.775 28.810 ;
        RECT 128.930 28.460 129.650 29.180 ;
        RECT 68.255 27.390 68.575 27.710 ;
        RECT 68.655 27.390 68.975 27.710 ;
        RECT 69.055 27.390 69.375 27.710 ;
        RECT 69.455 27.390 69.775 27.710 ;
        RECT 69.855 27.390 70.175 27.710 ;
        RECT 92.255 27.390 92.575 27.710 ;
        RECT 92.655 27.390 92.975 27.710 ;
        RECT 93.055 27.390 93.375 27.710 ;
        RECT 93.455 27.390 93.775 27.710 ;
        RECT 93.855 27.390 94.175 27.710 ;
        RECT 116.255 27.390 116.575 27.710 ;
        RECT 116.655 27.390 116.975 27.710 ;
        RECT 117.055 27.390 117.375 27.710 ;
        RECT 117.455 27.390 117.775 27.710 ;
        RECT 117.855 27.390 118.175 27.710 ;
        RECT 128.930 26.885 129.650 27.605 ;
        RECT -12.925 24.900 -12.605 25.220 ;
        RECT -12.525 24.900 -12.205 25.220 ;
        RECT -12.125 24.900 -11.805 25.220 ;
        RECT 68.255 24.650 68.575 24.970 ;
        RECT 68.655 24.650 68.975 24.970 ;
        RECT 69.055 24.650 69.375 24.970 ;
        RECT 69.455 24.650 69.775 24.970 ;
        RECT 69.855 24.650 70.175 24.970 ;
        RECT 92.255 24.650 92.575 24.970 ;
        RECT 92.655 24.650 92.975 24.970 ;
        RECT 93.055 24.650 93.375 24.970 ;
        RECT 93.455 24.650 93.775 24.970 ;
        RECT 93.855 24.650 94.175 24.970 ;
        RECT 116.255 24.650 116.575 24.970 ;
        RECT 116.655 24.650 116.975 24.970 ;
        RECT 117.055 24.650 117.375 24.970 ;
        RECT 117.455 24.650 117.775 24.970 ;
        RECT 117.855 24.650 118.175 24.970 ;
        RECT 124.930 23.660 125.650 24.380 ;
        RECT 140.255 25.490 142.175 26.210 ;
        RECT -12.925 21.220 -12.605 21.540 ;
        RECT -12.525 21.220 -12.205 21.540 ;
        RECT -12.125 21.220 -11.805 21.540 ;
        RECT 80.255 20.300 82.175 21.020 ;
        RECT 92.255 20.205 92.575 20.525 ;
        RECT 92.655 20.205 92.975 20.525 ;
        RECT 93.055 20.205 93.375 20.525 ;
        RECT 93.455 20.205 93.775 20.525 ;
        RECT 93.855 20.205 94.175 20.525 ;
        RECT 116.255 20.205 116.575 20.525 ;
        RECT 116.655 20.205 116.975 20.525 ;
        RECT 117.055 20.205 117.375 20.525 ;
        RECT 117.455 20.205 117.775 20.525 ;
        RECT 117.855 20.205 118.175 20.525 ;
        RECT 128.255 20.320 130.175 21.040 ;
        RECT -12.925 17.540 -12.605 17.860 ;
        RECT -12.525 17.540 -12.205 17.860 ;
        RECT -12.125 17.540 -11.805 17.860 ;
        RECT 68.255 16.495 68.575 16.815 ;
        RECT 68.655 16.495 68.975 16.815 ;
        RECT 69.055 16.495 69.375 16.815 ;
        RECT 69.455 16.495 69.775 16.815 ;
        RECT 69.855 16.495 70.175 16.815 ;
        RECT 92.255 16.495 92.575 16.815 ;
        RECT 92.655 16.495 92.975 16.815 ;
        RECT 140.255 16.470 142.175 17.190 ;
        RECT 104.255 15.455 106.175 16.175 ;
        RECT -12.925 13.860 -12.605 14.180 ;
        RECT -12.525 13.860 -12.205 14.180 ;
        RECT -12.125 13.860 -11.805 14.180 ;
        RECT 56.255 11.880 58.175 12.600 ;
        RECT 80.255 11.880 82.175 12.600 ;
        RECT -12.925 10.180 -12.605 10.500 ;
        RECT -12.525 10.180 -12.205 10.500 ;
        RECT -12.125 10.180 -11.805 10.500 ;
        RECT 56.255 8.290 58.175 9.010 ;
        RECT 80.255 8.290 82.175 9.010 ;
        RECT 104.255 8.290 106.175 9.010 ;
        RECT 68.655 7.105 68.975 7.425 ;
        RECT 69.055 7.105 69.375 7.425 ;
        RECT 69.455 7.105 69.775 7.425 ;
        RECT -12.925 6.500 -12.605 6.820 ;
        RECT -12.525 6.500 -12.205 6.820 ;
        RECT -12.125 6.500 -11.805 6.820 ;
        RECT -12.925 2.820 -12.605 3.140 ;
        RECT -12.525 2.820 -12.205 3.140 ;
        RECT -12.125 2.820 -11.805 3.140 ;
        RECT -12.925 0.190 -11.805 1.310 ;
        RECT -12.925 -0.860 -12.605 -0.540 ;
        RECT -12.525 -0.860 -12.205 -0.540 ;
        RECT -12.125 -0.860 -11.805 -0.540 ;
        RECT -12.925 -4.540 -12.605 -4.220 ;
        RECT -12.525 -4.540 -12.205 -4.220 ;
        RECT -12.125 -4.540 -11.805 -4.220 ;
        RECT -12.925 -8.220 -12.605 -7.900 ;
        RECT -12.525 -8.220 -12.205 -7.900 ;
        RECT -12.125 -8.220 -11.805 -7.900 ;
        RECT -12.925 -11.900 -12.605 -11.580 ;
        RECT -12.525 -11.900 -12.205 -11.580 ;
        RECT -12.125 -11.900 -11.805 -11.580 ;
        RECT -12.925 -15.580 -12.605 -15.260 ;
        RECT -12.525 -15.580 -12.205 -15.260 ;
        RECT -12.125 -15.580 -11.805 -15.260 ;
        RECT -12.925 -19.260 -12.605 -18.940 ;
        RECT -12.525 -19.260 -12.205 -18.940 ;
        RECT -12.125 -19.260 -11.805 -18.940 ;
        RECT -12.925 -22.940 -12.605 -22.620 ;
        RECT -12.525 -22.940 -12.205 -22.620 ;
        RECT -12.125 -22.940 -11.805 -22.620 ;
        RECT -12.925 -26.620 -12.605 -26.300 ;
        RECT -12.525 -26.620 -12.205 -26.300 ;
        RECT -12.125 -26.620 -11.805 -26.300 ;
        RECT -12.925 -30.300 -12.605 -29.980 ;
        RECT -12.525 -30.300 -12.205 -29.980 ;
        RECT -12.125 -30.300 -11.805 -29.980 ;
        RECT -12.925 -33.980 -12.605 -33.660 ;
        RECT -12.525 -33.980 -12.205 -33.660 ;
        RECT -12.125 -33.980 -11.805 -33.660 ;
        RECT -12.925 -37.660 -12.605 -37.340 ;
        RECT -12.525 -37.660 -12.205 -37.340 ;
        RECT -12.125 -37.660 -11.805 -37.340 ;
        RECT -12.925 -41.340 -12.605 -41.020 ;
        RECT -12.525 -41.340 -12.205 -41.020 ;
        RECT -12.125 -41.340 -11.805 -41.020 ;
        RECT -12.925 -45.020 -12.605 -44.700 ;
        RECT -12.525 -45.020 -12.205 -44.700 ;
        RECT -12.125 -45.020 -11.805 -44.700 ;
        RECT 56.255 3.640 58.175 6.360 ;
        RECT 80.255 3.640 82.175 6.360 ;
        RECT 104.255 3.640 106.175 6.360 ;
        RECT 128.255 3.640 130.175 6.360 ;
        RECT 47.215 0.190 67.970 1.310 ;
        RECT 68.255 0.140 70.175 2.860 ;
        RECT 70.450 0.190 91.970 1.310 ;
        RECT 92.255 0.140 94.175 2.860 ;
        RECT 94.450 0.190 115.970 1.310 ;
        RECT 116.255 0.140 118.175 2.860 ;
        RECT 118.450 0.190 139.970 1.310 ;
        RECT 140.255 0.140 142.175 2.860 ;
        RECT 142.415 0.190 143.135 1.310 ;
        RECT 35.830 -47.810 38.550 -46.690 ;
        RECT 148.105 -47.810 150.825 -46.690 ;
      LAYER met4 ;
        RECT 203.895 107.565 207.300 108.165 ;
        RECT -18.005 98.510 -2.890 98.810 ;
        RECT -3.220 97.680 -2.890 98.510 ;
        RECT -18.005 94.835 -4.550 95.135 ;
        RECT -4.880 94.005 -4.550 94.835 ;
        RECT 0.905 93.530 22.715 104.135 ;
        RECT 26.200 93.530 48.010 104.135 ;
        RECT 50.000 93.530 71.810 104.135 ;
        RECT 73.800 93.530 95.610 104.135 ;
        RECT 97.600 93.530 119.410 104.135 ;
        RECT 121.400 93.530 143.210 104.135 ;
        RECT 145.200 93.530 167.010 104.135 ;
        RECT 170.800 93.530 192.610 104.135 ;
        RECT -1.290 92.930 22.875 93.530 ;
        RECT 26.130 92.930 169.205 93.530 ;
        RECT 170.605 92.930 194.805 93.530 ;
        RECT -1.290 91.600 -0.690 92.930 ;
        RECT 0.905 82.325 22.715 92.930 ;
        RECT 26.200 82.325 48.010 92.930 ;
        RECT 50.000 82.325 71.810 92.930 ;
        RECT 73.800 82.325 95.610 92.930 ;
        RECT 97.600 82.325 119.410 92.930 ;
        RECT 121.400 82.325 143.210 92.930 ;
        RECT 145.200 82.325 167.010 92.930 ;
        RECT 168.605 91.600 169.205 92.930 ;
        RECT 170.800 82.325 192.610 92.930 ;
        RECT 194.205 91.600 194.805 92.930 ;
        RECT 202.970 86.080 203.570 87.010 ;
        RECT 202.970 85.480 207.300 86.080 ;
        RECT 0.590 80.970 193.005 81.070 ;
        RECT 0.570 80.490 193.005 80.970 ;
        RECT 0.590 80.470 193.005 80.490 ;
        RECT 33.900 39.930 35.030 39.945 ;
        RECT -17.615 39.630 35.030 39.930 ;
        RECT 33.900 39.615 35.030 39.630 ;
        RECT 32.800 36.250 33.930 36.265 ;
        RECT -17.615 35.950 33.930 36.250 ;
        RECT 32.800 35.935 33.930 35.950 ;
        RECT -13.115 32.570 -11.615 32.585 ;
        RECT -17.615 32.270 -11.615 32.570 ;
        RECT -13.115 32.255 -11.615 32.270 ;
        RECT -13.115 28.890 -11.615 28.905 ;
        RECT -17.615 28.590 -11.615 28.890 ;
        RECT -13.115 28.575 -11.615 28.590 ;
        RECT -13.115 25.210 -11.615 25.225 ;
        RECT -17.615 24.910 -11.615 25.210 ;
        RECT -13.115 24.895 -11.615 24.910 ;
        RECT -13.115 21.530 -11.615 21.545 ;
        RECT -17.615 21.230 -11.615 21.530 ;
        RECT -13.115 21.215 -11.615 21.230 ;
        RECT -13.115 17.850 -11.615 17.865 ;
        RECT -17.615 17.550 -11.615 17.850 ;
        RECT -13.115 17.535 -11.615 17.550 ;
        RECT -13.115 14.170 -11.615 14.185 ;
        RECT -17.615 13.870 -11.615 14.170 ;
        RECT -13.115 13.855 -11.615 13.870 ;
        RECT -13.115 10.490 -11.615 10.505 ;
        RECT -17.615 10.190 -11.615 10.490 ;
        RECT -13.115 10.175 -11.615 10.190 ;
        RECT -13.115 6.810 -11.615 6.825 ;
        RECT -17.615 6.510 -11.615 6.810 ;
        RECT -13.115 6.495 -11.615 6.510 ;
        RECT -13.115 3.130 -11.615 3.145 ;
        RECT -17.615 2.830 -11.615 3.130 ;
        RECT -13.115 2.815 -11.615 2.830 ;
        RECT 44.215 1.500 46.215 80.470 ;
        RECT 56.215 3.500 58.215 78.725 ;
        RECT 68.215 1.500 70.215 80.470 ;
        RECT 80.215 3.500 82.215 78.725 ;
        RECT 92.215 1.500 94.215 80.470 ;
        RECT 104.215 3.500 106.215 78.725 ;
        RECT 116.215 1.500 118.215 80.470 ;
        RECT 124.790 22.350 125.790 38.210 ;
        RECT 128.215 3.500 130.215 78.725 ;
        RECT 140.215 1.500 142.215 80.470 ;
        RECT 199.550 63.400 207.300 64.000 ;
        RECT 199.550 62.870 200.150 63.400 ;
        RECT 200.650 41.320 207.300 41.920 ;
        RECT 200.650 40.790 201.250 41.320 ;
        RECT -13.115 0.000 -11.615 1.500 ;
        RECT 44.215 0.000 143.230 1.500 ;
        RECT -13.115 -0.550 -11.615 -0.535 ;
        RECT -17.615 -0.850 -11.615 -0.550 ;
        RECT -13.115 -0.865 -11.615 -0.850 ;
        RECT -13.115 -4.230 -11.615 -4.215 ;
        RECT -17.615 -4.530 -11.615 -4.230 ;
        RECT -13.115 -4.545 -11.615 -4.530 ;
        RECT -13.115 -7.910 -11.615 -7.895 ;
        RECT -17.615 -8.210 -11.615 -7.910 ;
        RECT -13.115 -8.225 -11.615 -8.210 ;
        RECT -13.115 -11.590 -11.615 -11.575 ;
        RECT -17.615 -11.890 -11.615 -11.590 ;
        RECT -13.115 -11.905 -11.615 -11.890 ;
        RECT -13.115 -15.270 -11.615 -15.255 ;
        RECT -17.615 -15.570 -11.615 -15.270 ;
        RECT -13.115 -15.585 -11.615 -15.570 ;
        RECT -13.115 -18.950 -11.615 -18.935 ;
        RECT -17.615 -19.250 -11.615 -18.950 ;
        RECT -13.115 -19.265 -11.615 -19.250 ;
        RECT -13.115 -22.630 -11.615 -22.615 ;
        RECT -17.615 -22.930 -11.615 -22.630 ;
        RECT -13.115 -22.945 -11.615 -22.930 ;
        RECT -13.115 -26.310 -11.615 -26.295 ;
        RECT -17.615 -26.610 -11.615 -26.310 ;
        RECT -13.115 -26.625 -11.615 -26.610 ;
        RECT -13.115 -29.990 -11.615 -29.975 ;
        RECT -17.615 -30.290 -11.615 -29.990 ;
        RECT -13.115 -30.305 -11.615 -30.290 ;
        RECT -13.115 -33.670 -11.615 -33.655 ;
        RECT -17.615 -33.970 -11.615 -33.670 ;
        RECT -13.115 -33.985 -11.615 -33.970 ;
        RECT -13.115 -37.350 -11.615 -37.335 ;
        RECT -17.615 -37.650 -11.615 -37.350 ;
        RECT -13.115 -37.665 -11.615 -37.650 ;
        RECT -13.115 -41.030 -11.615 -41.015 ;
        RECT -17.615 -41.330 -11.615 -41.030 ;
        RECT -13.115 -41.345 -11.615 -41.330 ;
        RECT -13.115 -44.710 -11.615 -44.695 ;
        RECT -17.615 -45.010 -11.615 -44.710 ;
        RECT -13.115 -45.025 -11.615 -45.010 ;
        RECT 35.690 -48.000 38.690 -46.500 ;
        RECT 147.965 -48.000 150.965 -46.500 ;
  END
END System
END LIBRARY

